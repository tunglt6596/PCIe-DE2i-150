��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X������]u�.���\�KI�?�5Z�>�%i�v!����wkhO�������X{�ٸ��Tb� )C(���B��r��q��T}��4�I�����#U����3�;e,�y��R��=�TS�7W�8���[�) ���9��!{�3iDS�2������D�)�}#�z���w�z�����?���w� F���`�B����EZ�Z��y�x�D -lI���M������kM8�9�������%fK�妨i-��X�@��Km`�@��}��@�l�W�,����z�1.��er;�l����G $([{�4��dg�3�@C'hM�J�����a:$��L>�h��&h1H���(�A�|��33�_?�#��U8���ܚ�J��bvң(Kϸw��Ћ��c�u'|&�/:��qI�Y�f�,*�'�Z��Ԉ��|8�F[�}��:��S��	���|��òX;��$3���ZF��3��:�o�y��_����O�}I��-��fƮ�`����eq^��%%�#�?�J.Ŝi�S��D�2�Er�l�V���8mZ���a����%K����=�Q��J�{v�e���s�ƭ^Z^�'�A����W�a B��+�����2o��Ov
;T����%*H2G���utl�����#_xvt;��WD=P�=�I��:�� =�T*�*��+�#e�_������>,�t������ku~~4��&o�+{�6�:5���^���1x>o.�����*�5f	\�0���ӛ�کS�k�3�x�k3��! !�Y��:!��*�A��Nh�v_-���
_��x���N�"�Խ��A�-zP����V�Q?��p�ͱ���z�G�oZf�F<�l v��>ܲ������~�7l*tT��4�1y�WدWFqV�T�y���P�=u�6�B�&I�0Q����NF�,�U�����>�[ѩg�"80�k&��Ä�@*�ݾ�V�盾�i�	��.��8Ghlʕ�`�JW$a��Z�G�r��7�
����f���P�mi������|�ݡ��Z�f�$��zd�l�<y�U��|�h�?�T��iZ��3���L��YX;(�'��}2�
p�_�pn>�?�'t1b*8 A.�W���я)r�%e�n)�j��
Q�H���=D��D-z3��I�A��QS/�J�B�֡��z�rV�#���go`������=.��k��'~d}(TD\(5����տeH��� 7]Uj�l�EO�_�}�ҁӗ[� V��*�gWF��%�e�&'�s��ҫ���q���47���-(��ă(�	$�e�T�E� ��#�;J�",'_r�q���$yM�{�'�HF�x�.�S�d��M�[L�����L�=_����$��ɐC�����f��h�%��=Un��qҶUv�rt�JU�8(Mb�DG���E㽛�����
9W��Mrx#�DW���G)�_ǟ�jwGpi�[��̲F��vѬ_�^���-P�vIO�S�W��пt�	<���d!ژ���!�+u)g`�-��ձU�FY�.b	���.6�Қ������xL���	2�toܙOh�r"u0`��e$�nfa��w��6�R�ߤ�=5��A��%���2&$F�%�oO�UN��h�7{<������o`@AD�D��6�d�^N�U�]�qFr݉y��AjD���/�/���b�f>��֛��(-�#2#ӹ�O�>��;w�\,�\�,L}-���a��}�c!~2���"��ؖ"I��$	�Bn�2u�1�(s���xaf27k1�6+N�_[�e����r�a�I��ԉ��f�ޟ�����.�<��Wvw�Cb������g�� ���C�I�w2T��.�$pZ-�7;oN��m�b��>p0B+��f�9V�����G�U�(^Z
�\c_�>ܺ�l߬r�R�� /�?ީ`��x�l�]�ڈ(sK���Ćh�r�Uq�g��lϳL�4�'ki��C��E�!�fYit�C�~��!`�{�TP����H��t}mv���  h��x�6B? �{RnR��%�2������oL���#��vz@�{3��V
�?9P)?�]5�J���E�����2�_P�����{E�ӡ�}3x+ZC!�(����B����~���s���w������/_�W�H�y\|�p��p�
�^i� S�s{�PgpWV��q�'��'��%�!�C�y�r�㍔d��fJ)<��uQuX��,\ŤV�=��ŭ��)R�������T��a^��ɗ�+\P:�?H,j򠓪Ͽ.@=���3n�m�g���%G��V�X����=�D��_���i!cF��l=�YnIT��{���'چԚ_��|�� ��WaFFUJ���%f���8]�^nTe�̃�����{qY����)�36�䂚`�H`2�8Eī�vKr���S�yy&�j��c��F�߷l�U}%�+�f�^�� R�p/�ؼ�O�*����o��dm02�ʃ��Y�~��B�����GgB;u }9���)��� ��L��=Grm��q���g�%)�>���]mH��K�Pr��XVOW�s+~;t8-�X-����X4�0�[����l�ğ�� �2U)�؊�U��y���,��WLV���2X���\9��Ż[�̜�z<�oC����t��*h��Q����
2nR`�D�V���|-A�m@����M�9�>]#���M�����_��G��f!쒁�� �%[k��x5|~rc@	�[)��.L�OڃJ��h��RSkWFy��8?�ظ*0X�O��ե6�U�����4i�j�l���iH柫0���c�4$�����`�+�����o 4=�,�vK�-_|�.��*K�έ�b���ʏ��U��򴾿9B%���2�iY�-���}��w�^J�$�$�"��%~�{"�}����0�E�P:��1r�بQ�Y�f�%�s���3(��.w�.W
��p�RA��Y/�7!�����)˄٩�� 깢�E,�*<9r���4jw/ܚ�1+�j�W�S�#�Ej�4�S�^��S+O�^��n���N���5�ӳ�h�ғ7�0�i��
��G�1��'�[�T�̷�E�=A��>��\z�!�]�ҁ_�}�lm72��L� Nh�K}`��5�N�0�W)�}"�C�������o�7��<���*�b���� �2�ph��qǵ����w���aH���-El?c�A����*��v��������UO��q�.�"�/��(��i��y�!��Ezz���ש�dO
H �A�</m_��,��b*v]�d���H����1����7���t�]Ղۅ�.�?�7���Lڪ����^RQ(�+���������8��@��rG��6c�� `���gZ'
�W_8��u.@�]��-�b�͘�b����i�R�zvd�
�@�+ |�f��\;��[wY+t
M+������}D���;�*KG��p�h�|�K͋��7��>���m,����1��JW��g�!Ӽ�����	�BS{s�nW+B�6���B�ŷ��1�)�^x�%7���	�|�<� ;��BX~�^��c+FR|}��k�W���hg>6<~��C�/�fo�V�bC[\�|��[��SpB�C>M�e}��������[�"���<��c �%�rQ̾��JT�;��|���9��zY��k�JZt�M\��W�̛��G5���Fg�F��j��2�����!�ֺ*�'[n�y$M@�{��
ܸ��s�b�
���ʍ���G�cOne� �|�h����=��%̠����5�b-�i�}�o�|2l���LAy��j`���h�WwF!�Ƒ+���(�������t�y�u=H��LcS��K1M?�ڇL:�~l��z�%�~u
�+>!���1pz�O��B*|�X�p��M��̏"8ŕ�P�e��6�?��s	��rp3��D��Y6z�ռ�Y�����U�_�e�콖��>Z��3Z�b����ۼv�?L�E���oן)�I��WN�>?4�n�[\H롄�0u󊅘�ۡ�r�05�t (�5����=^�������^�r��16�:��)���AZg��/���ݗ��m��3a���~�i�_���`�v������j�;�|��c�(�)S�(I�7�5���ޓ�{�]+���*�1�)a#��I��*��ݸ#�T~Xh�.N���Լ�)و��f��x�ūN1ZΕ�Aw�f��$
�6����XP|�o��u�o^q��U�����tJڦ���Z��ey5;��Z�u�s�y�e��,uD��z����eu�����(eM���q���RC�,W������v����F}v��b\.�i�����v^'��mnC�%Y��zT�v2)��:l�����V�F�X���p��r��HQ�Ż�/�'�sHa��X���*�MQa*+���q�B�F�@XB� >С�}�;���B�kw�=&u��#Rin��k�:�_��-�f��`GfZٵ�{$5�z�п�n���s5৶ͩ�ow�kBk��w�9>Q�gř�b���6�ѥC�ªn��ZBe���bq\Ru��IF���$5w�ԷאYH/!��*�gk*��>X��3�Os*
�u��������F&�`�gD�^��f��*�_�Զ�m]O��$�K��o�`���X�vF=a�h�]d:ዂX��l��N��g�OB7QTV=6A�j�S5>�/��H9��T}����t0ހ�N>Wڠ.x�JJ�%��P���C+�Á.�<����8��L���Jn�@��"���Y��r)Yʸ��FSM����C�Y�R>:���1���/c������n�I�	�'^�?�6fW!��T�J-t�	`Y��Zy٪K��Z�
f����-�jD%r稁 ��#�FZ�yw%�ى�x�x�	/�T��ٹػݍ����ɧ������~�B�ۣ��~n���3�����ft�0�%�t��yZ4�Oܹ�������`q�,�8Cc�F� �2�
��3�ya��@`g����΅'�����,��w��-8�ځB{��<�4"ߟ[}0��(��0�=|8-%�����A��^�c;1s2k�2Nk���8�I�r��H_n,����MX��&�G�h �	T��)�)��q��Q�"D9��Vk���:��񽂷6���l@x	�R}OY��C���0J��,��;.�'��4����>�ֻ�P��o����#�ܱ�sN[K2��$��A.���>�zL��Ƣ�&��`��Pư�q��˞�å��T�����[����uߪL���*C����z��y�ΓhwH�����|�3�a���(��]�ĳ��;-ZǼYǃ�r�o xI�͗ �鲜̶�I��]�dt`+!h�'�\���F���a)"�d�{�$%Л
	�n�9;�DY�|�b�/·V��>���A L��%֛�g]#���s%|�r�d�lD�HLpg�['r[=�����V����0��&�6�mZ��y��v�1m{QS�~�8N����
}����UҔh���)�j]C�\(�73�~k[V���V|:R,�U8�|ƓȽ��~4�=�� ZO�HqG���k�s#biC������[���n|M���:�������TN3<�S��s,�v�@��>�[�9ʉJ�(��
XH���ժ]��<)cmJXG�je�rL�N~(��@�㱭3�T�V����T�����Q����H��G��'���=N�N��-e�W��yD6v:)+)�kY׏��)�v(��	�׎��s�Ce{ ��%�Сz�w��P$?)�ØV�v,I:b��3�e���g՟��g��SR��sF2 
�_�4?���eT��犘JZ���(�(���
�,�o��b�=rկl�+��;������wi�a|�#{C:U�{,�����b�0�3nv	���$��wD*r��|��81^���D�M�@�C��!�_$%�x;L�4�i�*�2a&ܫ�&"n�R*�ǣ�c��,㪇0��A(�Փ�o~�?c���b�����Y:`K��Tq�s^&k�T�=���e��6��W-	�t�./���t����TS������L�t�w;��o����;����ˍ�^Fh�Y
�g�|�ZD�{��$��qX�+��E2`�aH(.�^� J�Y�i��5�H�Q����K��,�`o����ʎ>�tE�:2��Mg�L�K@lS	^�����3������dP���M�΃����J�2�UGt��r��C6��J����&��>F*���׎r�8��K�m�������΍jT�QTS���Xf� ��J���[h�ih�;*�{�+���AtEkS���7�8\"I��G�V&� -	Js2�*�����-�D�I����ɂ�߾��0�#�족kY5��ԶI��po^�h�.�#�
@������-l��;�|w�f�J/1�w���|.�u-����7�x0{�Ԗ`
���D�O�k�Mb9���##�c�*�(�����~sK�mB3����W����Y;��'�Y_���%�{^fy~�t�K�n�)��A�q!<�%;'��R��
�)>�w\_gz!���>u�@'�m�fsH�Z±��׼��#��j���I�cU�_��*"��Kj՘�^�˭���~���0�%�I}��7�_8_�?��ů� ��u[��Q�\�Eq{;����K��I�G�J]�Y�K[�l�%������u�h�§E.$P��=А81�?� �N��'�a�eT�C�^����J����x�ٍY�s}ՙ9�V�Ҭ.���wv�i�FKO�.WXgNC!2��3��"�sa��b��L%��F�p��W��q�Q#�U�����w��t�)P�\���Q�o���p�Q&?Թ�%�c�4g��@�cLB�G7p>W~��WD>�N�����?W ���__=:;����Dx�A�Ǽ0�tU��+��x��~���#�WJMצK�� <�x� ��欪u��� "h�e��3�����{�q��{����r�@���SL*�)��KR�� }L�}x@���0fv�r?@� /)H��&�5�EK��>�l"U�z�."`c�;#�0�C�x�� �?�^E'�Z��g�gQ���,��1�m7���0��v�v!��.OO=����' ����R���u�oX�" �`hGW��r�����lt�U�q~X,D���Y}%�$����aJ�9KK%Ko_���B�W	%b5���0 t���t�XuԠ1:SXɘ����,���-�}A��@���NW��O�ߏ_P\���u)2e6������UÈetWR<�x��Am�[>�o���oߨ��-�.
@�nCX���5we��h����~���\� �\{�9��'�Q/�I�'��9JWy�h�����5�pL��g��5�@��4?�%5�p�U�Y�!E:�o����;�x\�yQ��>k�a�7r�zp�b7�X|2��ݍT�!��b"���I�uEv��#,��Ȅti�1k@�:&��9?��,�8����+� tX�rcGP�U�FB�l�6�
���YS_&���)N�Nn��h�	�(��@��iP���Nw�JH��4�PCЯKꎽ�W������R���8�����Aݤ̰�Pq$�Pѣx�T �g�i�|=��}O�;��w���=@��E~�8��֥�HZBcn~D�R	��?N[C����CeF�� ����h�޼p?{�'ė�����*�X����A7����{q���:	z�̂�K�ِ�YN*n[��
Eb�!J�c�ό���WI,�����-�k��Ua�:Hf��{2X��T?�u	[�;$�͏ƀ1�x�%�S�j�A�ⰸ�Ry�b�4��E��إ���v&@ɡL�C��,��Ǆ���m���X�cGd����.����E��K��
#��P����$,DЎ_I۲����R@��ii|�oZe����|�!�m�ʺv7�_T�I��v������up��/��_3H!y�w�@mÍ��Dݔ�|J����(ҷ.�x!#ӯ�R��{'��'�"�&�G�*�W�^���Ң�8�������1����h��;��u�WU	ʳ}�j'>��ŗGq��fGpS�B�����f�D$����*���R�g"�=ԗ�ID�{,�q��/i�잷�s�)y	��?�G�~[��˝�g�� f臙����lϡd8�O�>9��/��������pɟ���FW,8f������|Z���m�B���V�����)-��'86U�&/��^c��V�]ЃT��3N5�*tK�Z��(Q>���B!>��GNV��$�;�z8�Q��ܺuj�4<�;!؊�Q�"�����J�D�;A��m���;+C<[���t����h�kn��Ґ�̈́�Ɠ Rm�d��Hбr fp_��>]*�T��[��v��|:H����.�ޡ�����A�_xJY/�f�x,�QRT*��5�- �4h%6l�I:'��:Ba�W����mK����:�E���>ܞ�S͜.g���;{��K<6��wbo%�}�M=�v�{���t��;��q��#9�� �֏�]���.�7�m��LS�4�p�0�R��Uk���߭kOF�Ѭ�P�5d;�$J�3��]Ng7I�i��l>;Ξ`�V���Q��,ӁZ�A�9���
�|�)α�҆�xbQP0$���ؤ����#�f�� �}=]/ɠn+ı�k���F�2���)�8ǿ�Y`	Uͽ=�Q�ωKI��9g-�Ms��"I­| ,k�f(�r�J�LtFJ:��Ь��yH�Zp/a+���{7�~�c�qXϐ[Ȟ�4/ *���*iw��(�w�"���k�{e?�ת]i����/�O�<8�Ð̀�~��!P��6RF���r�p�l�:�Ne�E�B��eT0�w	��E�k{��K<䶨�O#
�(���~bn��r�]�؎���gSIL�x����`�BjN��������^e��}����A��?֜@Jd�Y���vy��	)}	�xK�
�]�eH.ܰ���9J�I�O]
���d%��+�r���G�ʴ:뉊f�$��|����l�x�!�\]5�W��u�K3�mY��R���+O:�G��އ,�(k����d�-O�"h&��(kf�y&���8W�I����v8H� *��C�.�����5}�&�2h8�k ����u�������\D�Z-TM;>��*Tƀ�Y�J���ax�Ԋ�'�Di/��c����F~D�gJ�<��9��f�P}��e����/jA2�� �f����������2�6�o��D�xiW"��*G�����d;qM��j�܉y_�jh5�ѱ����g#��5��D�+׭�)6��;�"0�v� ��O�uɛ9"��b�ܗ��ꍟ�7���myp$�[�_66��]��^G$��LR2r5`��̓����q|�3�8��ET�A�@�
��m�n��ރ���]���-pjI�+ؔ,�rh�ȫ�Ek,��옭0\3�D�-�	����
��X���C�*;K�X�sk��"�!63�^���%�%^�e5y`A��i��0V3+��\�X>g�D��6.?�O�"_CL'F�ǘ`�W����>p>�l�qf�".�|W0?2.��g�(N��O�D�![j���r�8�ǟIi]8����H�K-M4��J^"�
�	
bj�\k�F�\��Z���}�:w �o�>��b�������L
��?M�zD�v�^��cq`���8��U�5'�Af�, L̵q�{x"�[D�b¡��`���*H(/@�o$�u����$��W�
O#j�R�s�|=�e�b� �g^��P�3�G�(��ڀQ�؉%4Ц,}��[��Y?�4{���(4L���j�7IIMd��_�P���n���f�W���z��fD���i��m������!8B�_#��Vߋ���ﵩ���L�ȇz���{���M��o�ԡ�o���	�O�}N�"p�7�D�K��� ����]IH�;��&����j���q�J����G9Y���py�4K'�a^M�kUUd2�&~��ϝ��(Y�b����s����}d���� ��H�jt9+N�<Ł�ס@�Q����$�Bu[��H��x ��x}{�
Ղg����hY���/֨�����Q�/�_�٪g��K�Βr�<��}��Ft;Q
L����c}� �)�o�@Վ(h��)�횾>�(���J���2�]iX����z�tN3��MD�{��S��=���	��HeM�(�m��"�^y�ہ����S\���؜����չ���@����_�l��`�! ��)>y�W0Lf�Å��&�K��#+|$�1H.7&v����S�j �o��V�0��;Aur�"��;R/���o�GHg���h�m"�է����c�N|�����U��i!F���C.�|��>��K/K���?N����˲GR4�A$��@9Dʛ�pk�#B�l���`e�}�^��N|�,FK��K����O����r)���4Aw�D5�.��\���Te�b�G�DU2iկ�9T��U9M�A�3��z���+{-�V��y�`kݜOR#���q`��$�.��O��o؆�i�8R8��)�"���5�RX��$���� }�=$؍�Άz����8�7U�c���۷)u���Wgb��-��I�=Od�ڛT���L�+�o�]Ua�O��n�eOR	�!}K�&^��x����L �@�Rs�&MW�z�D�b�'T&7'�S��Y~.��ڇ�w�14�(i��ñc��]S*_����M�#{��o���m�3�ݷ���/+F��2b;��0��@��eV�PpЕ*�e���\�@��\�=���U�'�:X����^�]m�x.���Խ�A�+��;C-��gf����`'0�mZ�3ߤ_P
�� � 8�<}��\C؛��{Q�)��`���c��>>�bǙ��B��ěքV��&����>Nb��%�C�oG�����!2�%��1� �6��  �:9��Ê�G�ҒIb��Q3J#��nV^i^4�Z��I����B�쫝�������h�x�@�?tT���!~���T�/s�@�+o� �犢�}>?ѕ���K9���K�r��Ċh�!0 �JzXXR��z!v|�#7���4�!;�ʶ]t���+�i;���W�MV���H���C�Y��9��KQ �˿a��K���kĄf��������_M`ueDAi�^H���7�@r�i�f�;�M^Ǩ��(��lm7�E��g����9�Yj���P`�W��6�A¿%O���Vϖo_�r��X�w<BԜ|4��8����N�+��c��:M�c��D��9 Ò��M�>��>��(�*5��ս��� hߠ�%��8n���NuP�9�/�fG���;�T*�3�Ő�{�Þ�VX#���(
	�c��c��$�� �8 '���>�����Jb�G@��h��O�l����Ű����)-�
��0,����A�02@U�G�
�n$N���[�9��ט����%���K�n�;}��=��QR�	�7����Qy_�Nd+_�^��-�9�D᜸&7+�l<�-<��f�s�'R^n@/x�E:s,���:{R�f�?��6��2�B��}3Rd�$m"a�+Nh0~B�Z�w�}U��EU	5��'(ͩU�t����K��W����I;W�d`T�d}q��
���p�	\a��^�>�E~XI;4�6��wz�<�ϫ*L�f���붡����T�*?Ā���ׯӣ�-�3L�uwQ�x�\���3o�C��ZU��:���T�����<4z���ۼ#��a�7���/�}`"ɽ��j�K���$Z%���7��S�`ѵ��w��[Oq�M�f�]���g����� ��n��wS�0�e�L��?�����3g�!+E��Ȉ4H�o�&�w~o�A���vQxd�a���8�0�<�����g�y�\2W���zߔ!�E,�"�a[��i��TF�^$^,n٦&V�#�a��4a���Q]�w�#g�i\'|�Gȋ�>
����������R�Sw�@�)�u�e{���q�I�d�S<a()���>�C���	��&�$�t4n�5'��#"z�� *h0�sP��b ��DC�`�X$��/k�J�Ⱥ���e1@i�2�u̾$���o���;2�hV�'d��Fź�K!�~�R�U�:�⦥*�dFԏwa��f`|W�x�넽����,/���at͓J��.���A�~1��5�Z��s�	�=�|ך�b�E:+��t�h�:�ڧ�{j�FB�HQ ��("�$#����	n?��ξ�����7po�4�b�^�pW^�Ӿ�����,1����&~��q!�Y�*�;Gy�3�Q��mh�$9��J�6�(�,�I�Unw�~�x���`��l�� b��"�� {�B8��?�8�r�M��B��
�d�8�`*��N*cxZk(�R�w��C:	�cĐ_*r�h��]a��Ca���|U2b�i���?CPǵ�:@d?���l���M�����ˆ�ThU7�������	�h�l������.�c�0��t>i��z󽪏.U��"��K��+)�~~�$�n;�H
+��f��G����0S�]t)84�:)
.(a�#��UB��zp��rć��)j�eN6�e�<��]�]+��b��:�$g�z5��X�[�!�L�	�S�;SCC`	[��ꬋ�Λ^�;m�q�:�:ď �{7��ױE�����0jo��#�=�����ȹ5!]�a����L<����0����GT��|��DN�EE4=����]"FT^'XB��l����d勶I?��8���@7P	g�J�*0���-%G�'�v�~g9QE�@h��?>�j��̇���4o�.�ެ���w�>6���e�3�>�'<�5�E=5��s@�k��I���ă�lT�$��;��l�mr��H2n�Y���3֑y\X<�#�F�p<{���Y/�Br-���8$�{u�^��m����"ڼ�2�>�6���/�s�0��-�1w  �ข3�y�7	���G=h������T��"�tR�. ��`�ĘZ�v�(�܆�[�ا��Z�9��n�<	�j�%�%�b�@���������Y�����U�:�Ml��ųd�^�o�1>������^ Ȇ���~��UW��d?��,��L����+OID9��'���o^�a�^��y��Ҁ�����mE'F����u:I�S�Ec�-M@���D��gHa*/7��+jU��(�v-���K�YY���fM��wO��?݆��2���>��Of8�TKZ�v)��n�w��˘��MR�fr Ċiq�����r,�J�D|��hl�O���e����Lp�?A58�i�ֈ�S����P+������l4�`�%�v���65o��zn��̮�������|ڴ�a.,��d�A2�@�Њ���;m��WU��	@ΥJwx�z�cS�P<��m��Ln�=�v �0҆Ф���뜃q�,_������Z!�PT#�Sǌӂ���If�z@����e}$� �7��e������"�I�8���k|}O�|
;��@ԕu]m=�� `��!��ƨ�1ϴYׯ{�|��2�w�!o��ؖ�iI ��D�e�����'����:���jj�F�Bb����T�٤U�� +����G��#��-ݷ!�F	N�VQ�P<�ѳ�JK�8ڭ�=��"3��Ȳkaw�� ������\�*~���?�+��A����wq��b�/��S�/�6!	�9��VV�+�o�"7�8��,�#F9��m1���>�W�25�i-���HL�A��C�B�&]��#1�ƥ��q�"�Y�v��(���)�O�"Kg�*�1��0%z[<+SQ�:�Z�^���<�Y�90{�"
H��A8�%�)��Rhx��l?���Ϳɸ�������SKWګ�a���b{`��Цgᬉ�
�G��*�����k�ƺ�~g�����"Y ��u�#�,��"Ux~\)��Dk���s��.-��ڭ6+�,��������R��Mm_���-(�����EcP���ߟ�Ac�x#�a
HKY��d&��-�8AK�	1:>��_bb��ʘpP;)�q3�r�E&4�2θ�R-򇗍��5gF�*p�| ��"\�]�2�t�r:�7ש�A�.c�$	����~�o�HZ�Y�R�����R�|����sz�JE;j��� �֘u4����)���rY�Wc�7-���e_���&m��4���K!��VӔu�e��]��� 6H������j��Z(�Su���$�v:�c\�E�}!�8J���<�UBR� ��*�.��:l�:w�<:%������s}�"1��TM�B���|��d�HWI��nh.�w��y]D���iG�^��N�k¸��>�s,|�6.J�Yy��u+<2�<��э<�XJ�,���
�� ���%��aC��ħ�gJ��q�^*^������)oN�jxJ	d7w_u�
�j����w�{m:1�Ri�B�����e$�xC��x�A���b��ՈA,&[�j
!�Q�no�_�ZO�k�hJd��5�R�����ڃ�M���$zh����]�0R���`
kv��uhϟb#��)�N�ٌ�mn�&	)�i�w��a VK}>��B��wPz���ñ�c2�N��AԑfA=x�j 7��jc F��~��L�o�yL3���_��>�WOQ��X58���c!b:ܫl�f�7�ο�!]�j��S�龑9����tH@>���V㽠W�b��:`�J푢��R��/�ݲ�CT,�w[�ٶ��m�O�!d�.	!�O�d�2�+[;Ɇ��!t�;�q�ҟ�OųV���g��KH�Iy����`z,Cn*Q"�u�5��?��hq�3�D|��$i�	K��.�D�9���m5����a&R��C=/NK���������Pm¤'�e�ßR�����#������A���?w6�BWD? -~�V,�/��"��dti�D����R�d�H㸏s�I�HX�np��Z< �����^�%RW	Jo�7����v�P��k?H �i��57J��H&p��"d;f�r��P�J��{-! \@f�⿳n���7����"��u�ח��ı�V���
p`/Z�1 �x�ݦL	<>��72@�(�[�#lo�� �x������~��f6�_�W������qe9�%�.5o�����[�o������|8�^�\t��;�:�׫�p�~Ov�+�W�P:����0�Z�h�b�zT�q�۪�芐}^�;��bJ|÷���T��$��`&�sc��g�p� ��:�('(�ƄF|a��_�+���bDh��x�ߐ�B�=��[���Y8�zk�w���V�Ė���|@�l���|���|�h!p���ßL�Ʉ���K��Tq7�j�c�&����� ��� �r?	�3<i���|��=|م@E��@[C �m���ڎ�QJJ��@��`��;�a&�ꄏL�a����1�Ǻ���0+	�$*�{�`�W�M�4�}� T�0�2[��y�le��-���jH:.��;��ԅ���hX���GXK�e�8�(�����f��g5�a�eF�G�(�����\~��HPb����F=N���v7C�(�=��ӿ쏢]��c�[A�W��Si�D٥�R�Z���]�ǘ�� ޠ�7{ϷҤC������cfl�����h��9�c�g�_���,��܌��|��S(8"|qI���[tFk	5H�|
�mO"Z��D�k�8��U��
�pN7�HQ����e��Ox�	�«�mP�A��B9����]`�oh�,��pf���L���VX�7P�h�t�!vᙒ�[���$�w��tU$� ;\��s�ˡ<b&dV3Ő�"K� ��"���2����ǯm� ���+ٻ.���z�*���9�۫�u���x&*�O��ܪ��{
QA.{��c���~��v�;}̻� j ���^�RX��ǵ��vk�$C�+"$D�� �I)��[j��zTcƞh'a��Y{3ҿ���4ϋ��yZ��ԿV�����WKy.@P�g����쐤m���M��lDXG�H��5�]���^����h�N�� #���B��Qq�u�#��`��f�6[��'����Z�Y!�i�T�n�4���r)�tt�"S3i�KJ/�$�I�[�%�t<b���~��1rK�x�L��'��h`wW��E#�����J�ۥl� T ��B��wL�^r`�(xqq?�z��X�`ͦ�,D�Nړy&���F)�Z�d��G�A暭ܨ�?�?��@ar���y~�Q���>G�ľ������c�Ҙ�$1�۞�FT1Vp5v�
�y�����l�$�Ɲv�Me�\�]�!G��Fd�S���M�B�Y���d�ӎ�17VeM��;����l��*[5��J���߭=�)u��CLkj��+}����8n�����5�g�q�L��Ho�4@�Y�.������>R�U	�'w
.�̻�"���y������B�4�%[�שJ�G}�UD���-��g��d�=$u�ݒy�:-'�g/�$���;��xt�܏�[t��)/GI������2�΂߅����e$�t���	S�	��+��u"tb�
[VݫF]�[��a��+��$�V��,Fn���7ʙ�9��)�S�������=����:Vu��y����&Ҡ�Bܛ˯G5���\�"�V_Ci�䁅I��
�%�	�E�k�{���l�ܖ�b�W�Y�0�o��G�$�a�_v��Ah��l����(F��){�����
'�o:ef�E�.�KZ
PG�Lv�֯QY�Q�PR�����4}w����Φ��{����qX���f}J��EV��(e-i���t�S3hĩ�Q�Fx_	t�ӄ���S;��4q'��8��,�i�(ю�le�
���Xu\�p=���L�Q�F^8��\�2�އ��O������j;%C#_�޼�,���n��]H�sr�'�z*L׵�u
}g��)#CT�K��^�����#^����PW�M��I�j�z���g�+�����p�Ȍ=��x�h��O3$�uzQ��N3�T���f���L_��)�1l2�ՙ5b��N�J��%Rw`@�� ��u�F�y�J�ź�0Za^��Ga�x��cM�t��ɛN*&H9O�\�� V�䷘)O�x<Xh���Ym9Y���W_���9#^����mĺd�*��(�M�4��BA(�~�[�-O�ˇ=��,�f������̓�'{��H���`�r�O����d�ͼ��n����ۂ���w9X9j�*�Ȯ>�浃K*sRRf��N�Vr�Z�Z��Q$��}�m�׌����!3�v��ڂ��DțuJ�O	�O��v�ģc����wN��Ғ%H�� ���ڛ��UpC�!յk�d�7���_�s&��"f;�\�,�>H���_dC�7��]����'�d}>�^��r@��R��A5�r~x1�R|n��:�.��wnI�2��qJ`TGּ���ĭ|%�Q�[�F��o&��Fe��9gx<�*>֎�:����n楀h��H��rD�*�x,/3�	�9]N���t��~�Sb�>��X�Ĳ7��G̵Y5�OEr;��I�g'�y)��l��~�K6�5~�Og�&���fN�_;@J��&�[�����㰤p���G*�ЪlEDT3�-�u�a��G9�ɒNX&u�*e8�W�Y4�J�Lq��%�#�n�����I�\�A�{��O�ŗ��F,�!u��,h��ӭ}l��6�2����13z���}�:E��>K���D�h�����k;�{��+���������Q�h�$m�"5y�ƌl^�D���	`�����C6�ۗ�B�p<�+#+�6;R=[l�����+H1t����㖈�P�� _镰�ط`x��t0n���Ks`j�����ci���	�a�;�l��Z���Qa,�]�ރ��x���c�Hz�}~j|��)�Y�2��՜ńV��ڎ��.d ,e�)W
��1�gW�Yj��=�+���(�σ�kq����}�|x���V%���o�0�0�t���uK�W��7�:�M��5.�)��������g��mq�!�1�0ā��`V������~F��pf�5�e��eA��J�]��h=ՠ)c�<��6�]�1&��<'�.�;��,m&���5��Ղ�8��� �Ä	�	p�3�n�)�W�����Ҏ�`��Lz΋(پ�1�	��d�:΢�s�rO;�S}���
�r����T��N�� �h:q���6G�1�U�2wF!4d�F�O��"��b���Y��f�ò'Ά�j���U-�#�bN����4?�j��k�\W�PK1\��ϿGr:�_z6��cX/���,�;��«�+/��(�C��S�_�
K5��6��6�ō闔"b��P��^y'}���w����]E&�&#��ֽu9{���V��3K����!V��H��b��y|1���&u�p�3���RVvp�gڄ|t+��V��@�������}������c�x4���ث��B��Я���4}�Y{=�"��G��ځ����( �����^:�3c�H��ћ�T͢ZX��������<���X�\��~Bt��pcu�2���(Jl>V[�^��'�2گd88;�W���L��S���]1���I�M�\7d �P���E�OL��� 3�IaG�)s�Q«B�]�P\V�ڌ͔7~p8(&ʙ@-(�x��f�f����&��n^�K���T��>B�s�֯���$���������_� �#w�~u�����-�6'��$�g45X����g�r�ڛ1�;�_S~r�+��Z.��@���=�d��1wE$�M�ZI�����/���)
�:���͹>%��в�7-_C�8d>��x�p<���P��W8����et�'�����)����G��,����pm�j������܃�J0�Yx)(�>�Ψ�`I�4@.#��6���#>�0i�K�>�����-�(k�FO��ji��<�fuYݠQ��.}����v��	����3���5�����V�ͳo�K$���ʙ��p+ͯ{�uzX�O����=�򲆰s�p��w�/�K�t�%
��m^ �Ӯ��b�Bp��ݸ�r7�Lޤ9�Yy��3 ��NH�P���}���BJ����a�o�$N��ܳ��O4
l*��\ �ғ��*��@�U'�?������݋�4S�k��[y�9R��>��",��Q6F�&vP�%��5*�3��kȣv�a�g�{�eg��@cBL���`i'��SyS^�"�[)����wŨ惸ͷ:����5�_�_��;�i�H�-��w��4�#�(��h�&-��)�ֺ6��k]e�p76(�b��z�&FE�(����$g�e[?;��Wx�6jӞ�|1�^�f�z��#�?%e�LMG}^�b5"Rê� ��z���U�	a�t ����p�]Ɓ/�/q~e���9-q���s�f�׉��	=Kɲq��l&�]�v��gt��j����<��\0%w��x9l�лQ�$Ac�b���V];��X͋�z������$�H��.��RBɥ��dz0ֵ� wr�o���A��j'n�a�� �cԦ9H��Ꭸ��L?[G��U�Gs?��b_�E����]�=��w�O�}}E�yߔ�0�7n�H���Y�%�Q��[v�iUt1�<UBdf�P�Jt�{�h�6M�����P��Y�Xla��(�z��ɭ1��r�[�4ö\���"+QE��5��� Ң��~�h���*Ű�JF��U_R�%��������"8��µ�݅2���s�
�m;�o�_��|��$��05��#�U��Pn63��o��I�3?��K,�[>�A�rzj_�݉>�qn->��	IfR�0��*��XpB
����8h��s�𗸮дu�[���n!�7c)��^�t�#&�j
�m���*ET\���U� ��w_��ݶ[��@Zg��?�D���kL/��ٺR2��l]R)aa�SC�F��:�D��˻�=VJF�qZ�Xo=z��6ח����x�G�$�9�(�Y�i�Ξ�?��|�L�/�M'���fG�ιt���Ư����T����!�(s��5�h�]1�N�:H#/��-'��O���?"�)o��ه4�� ��0��7]x�w�>�nK�S��`}X�n<l����?���t�����<����Z;����g���>�[!<�.�+�-Y�+Z�b�e6!��"h`���̱���v���DY)��C������K?V��d=e�:>��W�^���dq ���'Sz��ns�~�q%��Ylڰ*��߅��\� a�'��-/��*��5��% "�izޘz���I�O�������<�C����������I�Ӳ:/����2 ������<B�.^�x7�+�j�<�Ӳ�N�Rtmb����d�^��Tn�/��Ŗ?D�N��n960�0� ���+f�s�(2+"���&�}
��/Y���p	CH�n3W��0�f���|� �5��W�]&z ��x�K�FQ��J~�U���_}l[��+mtZ��A�p�����~�Lr�=�فx�l�i.s]N�}i|�p�h!��5��7S qe���P�F�G�5%�Uzܼ<�M*E$K�$�$8�p�=�V�������8��1�тpp��Q-�����h��N�l�O���*�������d��8kVn��uu�Q�i��
7,C�%�ކ��H�)@��|���h�G%�w�J�`JC2.��?R�Ƥ9־�zM������� ���s-�<��?9�I���~N���)���l�c��6�fS�c�)D�qy�4k6M�8���y��G;$7���Y��.��w�y�*^?z ��I>�|;�&Z-K3^���n��gכ�I�)�E����f&
/qZC.A��*�op���&�c�f!c�@�~������ꐂ���7��*L��_ν���0�Y��xS�J!Jtt��6����Q�c�87��DbO<��L2�QB�����ris�[Xk/��%5ma�8G�r������:�O���=��,�V��Q�R��!~�B��U�ud�nr����O��R�������<K5���PL�����[ړ�7�8�z{�v����6ebFy=��o�^���2������>�n��t!e�爕1q��b45���lVo3;`W�V��n��_��~<���z�u��3cͥ1@�08�ѹ�@�v�n�bvc;���a�=�����zs˻�)��|��ǛJ"������l�T��o��K���َt������t�	�U(ڲxY���sQ�[�(l��Ss1f��2����k���.>Y+5�0����JYA�;c!A�A�����EL��m�ڛ��Y?W��򱌷����/sW̅�Û�+��~�'{�"{�G*��K�r��KN���w�"��t�zCϖ�/�&b�q�mJ��JT��c2w�O�}�����K3����B�:.��Ա��I,�`Q:��e�/Q"��8Y��!�ޣq�Q!X��W�h�Q�a�r��������g��yRA4���+q�bA�U�}��6'�*-2x�o�6�X,	�sfά$(��di��U�ZN,�Ew���qt�r|U���!̵'�5�f.���f]~m/�w9��g�x�k�Ի��\dL�	��M�����tC��v�XGQ+XHOV��Sr�n�X%�3��1�M�r�DT �gM	�BBßu�� ��-g��A���;5��0hS鰖a�_����"ſ�|�R�?E˗_��"��/����S���ђNz\í�JL��D$!�����^�j��
Z�ʋC�g�+��*v�-�os�2\�de��&>�B�s�_~S�1t����|�Yg�Oޢ���|h���n�]E2^��9�^JWD��(��P���@����%��<��rߒ^�r�nBI �"z���R�aR� ŧ��LeY�(A�4��%{c����ak�ys�8ך���J!�� ���ƨ'kr2��q2fI�߲�2q(IR�]n$Ykdf�_�� �r�8�JY+v�iꪎ��b
��MHa\j�A�ն���.�%�`>�j\
ERS[�������()?>9z��Dl�!�S�Br����ib�r�U�)_�B�D�d�?W�~���2��N�R|�ݵ@6>��{��ZzOIP�Q�~egL-aV�D�D"�����S����<?�Sᤱ����!�������ku?�Z��a��&��N��!@���G�2�ڰc�	wL��l(.w엾#[���2�r��� Y�G�}V�{^�q�zbZ1��F��� D"��g5<�c��a�K�/�� ��z�uh�2�Q5��	�g<�@�_E��K#+F���G��c�qy�q����`�N��Xȇ����L�J6�A
KA�3�/��nE���7�*,���l����z�
�a�ḩ����������g��$D�����&�+�;G����&������Kǩ�E0Ǹf��=*S����[�E���p��z�k�����bcx����B�����	��f�)\�q�ه?>I���_� EƲ�q`�>��iic�՗��G~�B�h}�U��x�r��?�j�sk���A#��U�U�T2�礸0H�;$�E�l�|�M�<�@����޺#A�\��Y��*#�B���绊���Q�K��_xnȡy���4�cZ2��i	�H:j�vZ�q\�Y_t���5W���R������܈���'/f U��[Z��,�ë�L��UhS�h�J8� ��}�Qr�s�+L�ĭ���
Sߍ���AbȔ����œ{[5�
	$W�^���l�(S��$Ƭ�*~@�_7��Ѵ)q:��*��(U���+جB&��G���UƦ�ڧ��4�<)�q I#o��0T���HH��m���}��]L?!��J��v	�"N�t��iAZ,���
�O��a���D���T)\��~t&ޥ
tJT���z�:xֳq�4(W
)��=�� 84��ON�mQQ��HW>˙#�X��������Ӕ�=�l}��s(����/�փͭ<�0��r
M��߫��±a����|/�V�W�_0����=و?w�<�4W�c
�!�ܴ�ѳ}1k\��nUe�Δ�ֆ~��@ݶ��J���z�� tę�i|=xSpf��دd����p��C��	1U���Ȳ�m��-?g��T<E����"b��w�e�y��f3�צ���|��Y�H-�����q_�����I88�~���$�t*ĐQ�9��������
Az�C���V��ߊ#T� ���y�����~��E�P�������k�<�z^��Ì/���<��vzde��@���?� Xu?ٳ/ǍL��0]��X���y�*�X!�?�9읡������I��,�,e�/'Dځ.�)T�Ss\�"�A8k�Y��F�IGE�O�D���M&�Z��X޲c'_��4�U�Y�	0(��@[�hc�(A��/b��l����q������֦�R�E\칮ڢ���3���#����c��
0����LE���`���*C�ŕ������]��� r��*��ޓ�ⶣ�Akڣ��u>4���
�¿�'I(��`)�۸*^�܆��:��#Я�Zb��-:�+���p��rh�[-�ڣ���g���*� �6�2;8�K�
�cC.d��4�exK֬m��������q|Jwvud�S�H>�.�W�擾�����,����3�%#4Ę��+0��v��a���o����VI�t:��;��ьw#�64P������^c�=R���
�,��ː�HM6�������
e�+�;xVۚ�/�z��L��D���� ��$�r܃9|pNU�P������ّ�Z 7l�f��$+�J[��`U�9��\9����O���;� :=�K�M�*퀜,�����wr&"I�����%�ь��@�]�=y�U�-e��v��_���ZesA��8��Z���k��κ�r�{h�k���I�|IS!m9᷋�N�n`�7�'���2n}�ݬ� �!ذ�r��ԱZ����_#3�ō���{�T�!���Um6󸘎���+شE2��A�!<�K]��e�M+�2�l8�v9��Dv'���X�bnζM�g�
p��q�L��-�E}���sn��y�0�/J���(�_j�$�c�HM@���n��lk�Q�Х����c���r�{��6|�s3�$y�.����)�+�tD�l�2ӯ��e��p"�T ��y�p����W��ee���M�h[�D��Xd:�ލ�E��l_8�+�\�*UJ�xqh��s[c/�
�4.���c[��O�v����z�# �u�=�nr�g�^�um4����.�Z������Fi��'�i�Ӆ��y�U����ҁ<�C?��sfS�i�x1�~?��w@��;sʊ��Q,O������h�1��b0����q�U��4�{O��E^e��-���\Ǌ��@������k�ke���W}�,����P�ZoA�t_j���g�5�۞�f�z1��%]r����w����Z��g`PF�E"ƨ���h��&��7pP�Ȉؽ�o^�>q ��K¿FN�.^8�VX=ĄT)�xi�R�{G��g������=~?���`.��Rn;�}?�a�[���,�L?�Pd�ɽ�s�^�����?�k_�������mn��7,�8���0BLU~�h�8 ��a����}!�Gů����v��2��,����������R�� �K�����b��\�ݓ%?�[�!�f^��J��n�K��W�m>/@׾���%�%�O�T��f��M�����N���'�G�(�|˷V���Kܶ���Q���[t�A���#�@��^�Ts1�LO7U���@Z(B��th�2�v&$�������jP������c `г3��\*�e��~�1��%7| 熢�O�g�o1kL�5�d�PA�\ὔ����	��"�i�I��sX,7e�ɑ5D���`�������2ɡm�:bf)��jwn|%��fyW�-�/��@]^�!��#�!��	�5���h֔�м����pI���;��1��#��)���C����*jdh��x9�6�@^�?J�ƽ..�f12��/�^��
PZv_Ju�َk�7�'`� ��8�MM�\�Ņ�cr�J�����D��D��[gmMۛ��b��_�y�	�u��D*��X3�Ϧ��k+�K3o�M�W
;	�Wҍ��rq/��2���pA�H�Kw�V�!	{��c �0$��R^,�|�2�[x��[�����٤�4�¿�p�;I�WNz�X+����8q;;��n#?�^+�b��k�c�V����uM��:��@k�&gݶ�,[�G�6��#U)���Ԕf��/�q��(ƭ\k��gN!��"D/�hEU���r�lUa�6P�nQ�JET���j���q7�"��g�2�h�vU.[� у^%�h������'�V�w�ɯ�����;��;K�:� ��+�X����k����>9L���ݤ�N͠N�m[�D���~�=2���u�͌(A�\�o��.� ����cԛ��>^U���p}��}��Y �i��8��#��\Bv�����Q�ZĜ&���2c��0q��B���S�t��XkMtH�euu��[�cP�X�>3��&a8�d9���Rg��iSR%�c�����C>���[1�ŹSOr����*�4{��?p���Te8�o	*�7:$47/�L�BD�>O���c�Md�ź�͘���ˇ�b���1G'?\���[��W�`u�-�����ۣ ���G���Sw��(�x��v�-�
K��L{�z��)G�G�V���~�g����A�߷P�L�Uj��S�ǐ�w6+��.�O��6-�"�k�A�~�5�f���ฤ�J}K�c�M�n��[��e_����|�#Q��q(ey���5��n~�s�Ts����/ٔ7ix����Ūhdew�n�cZYU0կ��B��$�[H�`�xbnU�)BQgBS��3dX�M��Ie[�	12A��U~�L��9�!��ӹ�f����l(Z"|;N��+!�}+�����v��ܕе� xDa�ۗ�j"2�,f���f�0M�<n��=�Q�K��*�yo@5��#@ (��d5�=�2e�ƁvOY�|sܤ��2#�b�T���T��}��' H�z��������>w/6��NQ9W����j��^�э���-��k#I�,`X"|3�+���i��'�>��*�D-B�汚�ѺC�����?N�8@���1J��pQP7%LO����\"G���Y?x�:���Ҩ�v���AsГ���S2���WrG9V"�p[���ό�'~�U�g`F!���`�H��	L�YB�N�,��+,�����Jn؃#�m���G�'%^��؏���(�N�g�$O����:ʚe�./mP�*Dg����QoW�Bd���l��hI�I�n�VJ'�d�iVý`C��d�Q2*�Hg�S��B����>9�t��5@��͗��0U����6:�n�j��q?=�Iy�_H�k~{6І�Z�:BM�)��`�*Y�.��:�b^������IasT���,N7���Qt�OX�b?��(E�G��<j	ٷ
�2��,��/��a�j�sG[��5��u���z�+d)\��7��RXu���&���u�fZe#�?�4�˯~����B��]ەP�oqpf��V��\ժȡ檅��:�J�x�[�����ֆA&�1��Ä���%�C��+�9���ޢ!���ek��AO��Zc��*��J9
�u(�dW��־g�ˤ��`E-�f�����̫%hm�p;*�H���.ru��H�������N�;pޅ
����3�Zx].TߡD��0#UXC_�� ,u����o��_���{�[J���=O�@�N�}��(Rz�]u-f��������_�D]����&���>�}�ʶc&ڌ�T�[�5c5���o#r"��:q��ಁ�5�Y}#�5h���������;Y�t�{�ED�D�q�7��@�)�a�ۇ��}G8�Z�x&���l�3�-�Pg�-����3G�v�H��hE�X4-ǲ�X�ѻ@��0p���\��r�90d�Z�h��@jž_~m7���j���py}�;� ��/��� �ś�bj���P������W>����rY|�zF�*N~4�A9k��{�	/4�
�R�>	�6: ��6�v"���|wojXҦ̽�i��C`r �i�Cٍ
�hۣX~h�ٍ��2�Ȗ 82��_�$�ܩĝ���|��������^e�a�ތ�Y:�$���C]F���\��=CQ4ф&H��.��<��b�u���d�m''���o<J5��#�hu������)S?n!b�Б2��8�7�>bd��Xv�$��[z넅D$4�f~w$c�$�(c��G�Q��[o���Æ�d�|��kA�Å�J8:Yr?�P�c����V���O ��*2ｒ����Se:e�_�����p&�a�L߃�A�&����<Qv��BO���Xm�x�m'��r��fGߒw1I�!1�d�'��~'_mw0�j��!.U?	A�����C�[����׿3�f:X�..���x�������Q�̕劢�vd ����m2�~�������;������d����n{������g� �P��j�h=L[���bܠ��:Q3�z{	���N;�M�K�_�_�	EVq����ސ�U�H�=� /���?-
���#)-�Y'��R�������_����h�j��FK�"���}I�/.��z�L^�svN�,�e^�U��(d/x� hZ����B5�j�'K.1Y�)
�}e��jأ��Č�ѧV��1�c�ZR0��^�>��N�t��D{��`�,�sU>A��� ��\^KԘ��[��w�N��9���z�N�DFH'k�B9nW��)!��6� �X��mP��B�=��@(�u�t��'ҽ�O��it�Oi�A/�w�:=Q�\��aX]%��;G�W�?8�i@������`��?Ba}��UTɚ%�kX��3OS���V�Z- @/�����x1�M���3�Vrw�9L���!XR�@c�G&��ѫ?�=�R2�ݲ���m+�`����d�ؚwc`C�妅���B>b�r��j׽f l�%I ݒ���|����xn�s���6�S�5R�ퟜ���r��MGY�(\y%T�f��-���cf�d3��yG.��<R�5s��_��$�}۠Q��~Gp�h?�[�p�ȒS��9�� a�M���rMốQb,
��.^p�$�|���P�d�M��ճ��8�	d@s�V�|�s���@lB�?��E��b'���v�	'm�Yt�ɷ�`+�Q�1�"�C�F?)��b��%!�->6a#"�8{�f�ԏ�A��)a@~qE8�+(�K��ȸ�ǌO�%��E�{,f��՝����0�5�H����p����-3rY�	� �n���~�-�0�.9%,ג��A� �m8���;����k���]���Њ=ź5x,�^������Q>��ݲ΃F�K�3�	������`ܩ��=��J�g6f�K���b���:MVk,oȽ�������t��*�8�ީ����T�nxi4�]���H��,Ga�OEp����7���-��=ʄҙ��=^���t�^�v�BO��Yu�ψ�$�z�sȆ��ؔR�E~��.�;z�y"12�1>�y'�_��+�xMA�K�	��ƟH��jA����6���=��Yk~���k��1��G�Ok='7)5�nm5ד�y�g;Ύ��AE����t�k��	����9��9�0
E�4�b6�AE�J*ոzP\�
0
�T�\wd����$�"o()���ْ{���y.���f�d�{t�2�*��Z�>�Bt�����jԚw��S��Ep�"b�j@����6-F�W��}�hܻ��9���lB��S�.x�)&nr;N��4	I*]��O��K���Lo�:>��}�׃�`� 5mV�����^��uω8�wlP܋a��'G~r��F�����G̈}�q������i\�A&��Ë6r��&M������/�d�M_�x|����D���O9A�P�j��$�AdF��m����v~�{���|������It�7�zL"	�09x��F�I%�Jrc�������!6�`����1��?�F1Lm���Q��b�����;�0�Ӵܒ������-M�7^�{�8���Q���|�;�g,!��ɣ��&Nɞq�K۝�S��`o'��g����PE+z�v>�߂����Puab�'�tp���5�3�&�tcݒt(#�5�P����	hl�=�Z㚨��D�z[�dKxXe�_/|�2�C3د�@>\���vD�����s�o�
٦ۮF����Y�+v��T� �H��'G(��C�B�m[�0(s��jC>6��7�T/8�¡!��'���s| �5!�����̡��!q��B����s38�`�����Ik �4�G�t'�f��%E���GG�F']Yc�A�S'�+�=�r�L�t����n���l�y7�GҢФ])^��Ye�vx�Gt�baG*�X�%c�z��@��`���jg���ه�E/ˁ-��v��/�~(*@��sui(� ����8p���m��W�(r˾H�$�0��7P:X��4T�jg�m���`���Ч
� <�=S��]J���r������
� ��ծ�m�_\J?᧫�
S��X�ml����o[?I����z

�أb� p�	�ǞyZ�?d&��`ޕlOЈ���n�G�Ꮾ�̳-+B�K/�����Ꟁ~Œi�H̷,��",(e�a�HLk�rtB�SExNeܨ��ϑ[x'�F عú�#旾��T!aE2{͟���� k𦱊�je�>J�lK��-˧r�p�y�eIpZ�:V��p#��dB7E��ZJe�8���&��}���U�%vk���2f��0�=θ��|�B�sD�R��U������Ը�ץQ�$Rx��� �F;r��L\e����E����6�J����0�J�$�}O=�*�����ҙ���?��$(DH�k2b ;�?@���krhN��ihQ�Z����Jhsf�)%�
�/9�e�����}Q�Y�T��{��f��1ތ�|�*���zTE���TL��F$1RQz��y[D�5H�e�����X��}<k}%�f�U�"�3z��v��>�,v�?S���a�U�t+",��U�rf��e�E��t��Zp�Fa��������[��s
b��.�s����i�!���Ay%j� ᦌ	�Pl4��@g~����$D~v �2 ���C�L*�gs�ƌ'�����T�%L-�M]ԩ�)� �z�܊u_���rk	��	a���������!Q�Z�� d��7�����[ÆQ���ljC�}BX��o��'O������ W�/�@�QC��9'� Ec��%l#��DjN�oq�6�d[��� �唚�^p�eV��@��v͘��9�T�;�*��q�[W�$G�	g|Dш'~����(������|�=�)�Z9XsJ[��/����Ⱦ��ZrY��,g��S�_�Q���UL ��
QS)���W�EЁ�L��zɚ�c����w�����6DH�2�	!��ҀUț�B��l� ��A.���~N��hX�[G��ů�+Ni�	0e��B>��lL:-ۥc�����3ԌB�󷎹�<�C����}̚Ò�x� �|�\Xt�H�3³�Eh��C�xȻ�aq�a��y�p�qA��8#^���I]�:�x�展O�P0z�#6Lc������9|��H	�D�W�j��J	��V'�s�ٵ��9�|��a���'(����EރM�gr^-�b�i�˷q<IxR��[}igNbs�]O����)j$۰���y�p�Z�ŉ �v\4efl'�i�zb����<s`�2�%S��nI+D���k"�Y{{���t�i�GR��햟���LMDB�Tܘ����:���>��{W�_�D��,�$��A�d�4z�9�O�)J�������O}�(H��()���T�!ˎ�C���Ӝ-����3�����k�G�)�e��ָ��OS�	�g�
�Gr9�JN��$�������No�c�kqzy6�;��	�eϗ�f@{�ԏ�����
��2�`[��c��?��	��PX޺N+���8
,v'��� �a��4δ�/ �!kI]X������fYv�3������F�VE�#2A����N���M<%�3��4��[�K�.'���0"̑yw=z�	��O뭩�^V
���E{ރ&��MFT�H�V��*u}�"!��с���'k�_8Ӥ��Qf�ǻ>7D��.�Q8O�,� .@%{�N�V�&Jl��%�x/�ؾ�'y�:���fs�&o�l��Py������d�3�R�ɔ��[���+Ya̞/�Ȅ0=E{!ji���{��s�+�>�N�C������!����"�),�=^4�$�^p2��(���q�����^%as�4�1���%N��e�uğ��*���A���Y��>��u�E���>������#8�Ӡ���W��Z�tQ^t�;�r�Э�f��3~k��]ݗV������f2�{���������[���]\���6�=���Kjc�j�b4�1Mk��E��~S�<�ɄP�2���!O#hL���� u/{���f�H�U"Kod��h儸�:Sػ�+�)�K[鑏��H�e�����I�W��j��"v�F�/r�u�U�m`���~������+�'Z'�5A�)ػ��@M�3��l�)NZ	����ur��ܪ��J��"w^	"�f
Qj�|+�,.5�u�5g�0[J�������! �N�y����h-t�,�(�lV�MT�1��=N �	�{�����Z��=f0 Y*���C��)i��[�]&K��K�L�OƼTE���� j��[���M��^O�~�S�������<�V@��������4@K�~l#;���Wd�#�81U0�`��40���Y��ұ�Zj�\w���V�3?�GWw�R��rp_8Z@,���(���`�IV�EG��o��%���3o�g'=S��\�. �F*���)[�����D��g!ڲ�a��R@������EG_����s�-?I"-��<�ʶ�/���q~T�B� �:�/n���ܹ�K��S�_�Ϧ�9+@���0�b+a�CF`���w>�q���2�&_ȤT6��ޓT�$�<w��(����:ѳ��n���}.�Yޓ�����j�	����Rڋ"U��r�	f�{�C��ߞ�O��"L`�h��v���px����e˜�
�a��Hъ�b�i/P�U�����Á�Z�[t�J��$���;���T��F���ђ�V��7H>��W��.xk�t��ͧ����Q��xs��n`�Ta�A�J� %�[[�-��,B��1�f/�O��ĮO�����N�^�{Ix�@_{�W)�f�:��.��NR�vE� �K��!�H�8$K�r��t>���-#�z�9�冃��uY,�q��y��>��:ܘX�Tr�[!.�0�X����Q�Q��cdfV������F�_�qk�xu����6�a��a� @'h�<dN�F�!� �u�*��k��>BX��fV+ƛ�;��!��Ι.�O�4ݫTi�5Y�Jn��Y���Y/�(�ͦ�9�(��Q#G�ӑ1)Y����z�<zYfl~_������<�����	��oN��"܄s��Ey�(�����h�"@�O�b�s�<E&�<��M�hrm[/�����o� x��>uw�f�r�ˮv~��`�4�ue�д=����i���B��3�
�K/z�7s]��U_R�����+���!���ff�]�9����Arn���?�Q��W%iv��s�v��;p����W��R���Q+A�EД�sF�.P�0�3����%$�5ڵ�'[��75�m�j�J�]i?<��?`�T�U"$�H�A�D����4C�{%y����6@,܏����yop�����ɣ�mfs�]`�ME�����|b�$1Aw!���kc�fϩ�x,|i� +i,;9��7�َ���p��ܨ�6{;�M��13!�'�:�������@�4���m*b4a8��h����Ty7�I,5�
���[[�Tt�9z��t�/'D��g���0&��]Æ	"�}L�k�}[E��Z��d�O?���G�E�����U)�u�v4���9P	$�;��
� ��X�kZb��`��׮�J5����8.O�Wax����+�~h��p���!NtIg���Y�D '*�p��g������o�L�����KϽ^� ñt�v�>n�l�W��n�3�c�C�J*z���9&�-0*\�=��������T���Ƚq�򫺣z	 .��֎��ۑ�.'������5��Νho�&��̷�c#8�G�`�E$T	oQ����!<�;�jx�N�q\p?t�O8U 6[,���L��B�M�D�`�y$��;��k����������~S����6�S#�:�z���VJ����|��6�L��fE��2�ۺ�~��d�"��}�p�����z9�Z���g�>��o�j��fh�����;�
S�K:¥b�V�L'UP�1ފ]��;�^��0�o}�*\�{4�겪z���mn<0.��E�s%�{�@�ϡ�2�����l7N��2q��c�d6<55��X�re��U�Ƭ:�q<X����Li<m�9Aխ.��T���\@�U��(��^"NR�D�2e��8L��\�q�( T����ǂ�n��$�l��5H��U'��w�AaID�s��$u
��h�v�Q�ORj��K� ү��G�f���d<WY&�h��N���f�7ߨ)h�Fc{(��[ض���W�j��+��8�
��g�ɀ[�=г1�2���+B�����{X�z@�$�?*��Ik�=���A���%X�D&�	�d�rt[>T��d+�k�/CLea {]��:A���V���&$	7s��.��3�,6�:ES�n-6@>1�t��%��N��",	��K�&%?�"����_�o���2��0���"�:w�([R���"���0V� ��C�Ķ{�2�P޼VTᤀ�Z^�����S5����x��u�&�1akOj��jIr��޶ޞ��S�6\hӎ�ɥ�!f8�q��t���n�;,�3� �J4]}ld�>�4�<�0�?tN,�6P`߁_��Lw�m��Ì�u�~�J#g#�M�oI��`����\���t����z�E�M��@�� t�&G0j@=V�� ��{�E�|b;.)��`?c�*v��d��+� ҕ���k`�g���Okc��(X Ƽ���zRF1�����Ȱ�h%�jZp[�=���W0����o'}|��0�lp�LC;3��z�>n��t�Զ~\����� 	]g��������v���,����E�Vў��Ub*Pq��Xԭ�*`��Z���#X��K�>�����Ƀ���p�Jff�R�/���g� "hr�J#�ދ�6.y8+�OQwX�\�J/ut3���H�+8�2�uŭ��~�!�Mn�n�����8���y������U���s!���P�k���i�{��3�����3b�z��M�����g�\̶2��eP�5 j#!�����m��z�����;�8�{-3IP�LGİ�Q�ܵF66���5r#���37��/��y �RY�m+A5����_C��~e���o֩�3�W��蕼�8��x>��<�93�����ӆ��eD�*5h��Ax��F�'��bxU�oW���mB�q�����k�����Qh<Em/�H��.�{�s�6�0��g�������
6��Vg���K�PXA��](�}�g,�u�E�5��&���(���1�� ?�g\�oj��Rz�jD�%.Z@�Z;3"�µDo5��~U�W��d���N��o�'�䩢�"��ň4U�J�X^�&�h��g�͗nh+�~���={?]��jlG��k���<H��_����(����y&h,�
bM�#e0qѼ�E����O�ͭ�ȢT'%M6)����j�rh�KԟTnϾd,�����vQ�ޖ�fI�B0�ѵ�@ߏ��.e�x��aș�kZ�9��0�l��U����BV���gUt�m�+Ea�]�o����>vT��CI��#5�ջ[��n���1�y4&��w�w+2�S_�K�_xL�P�S��ҵ䑟 �WY��0r���'�=��J��OA�zd[h1'�	��G%GQ�$]��O�O�>���-���uH����G)�5�#F��ƣ���Ysi�W��BP
���4t�l�v�������@�!OU����<�U���L�x���u)a*��%��XD��)+�< |9��/�q�������e����@�j���z�˞��F:C^�!r~	�77��^�3�Q�ͺ�S��1�� ��Hl��b��>uE\P(�,�cT��02��o��T(�s�'�T~%�#7�Q�1<�j�#�O��IoC��,T���Tk��s^X?��~8"�n�,����GᰠL�рY�
H���j��ڭ��ڔ$_-�dЍ�ce�rw���ʂ��=G8�m�{����T�Q�#�gte�<���WW�|L��D2�,���:3}1<�-n�a_��k��n�l�	?����}jiI��m�8?̻�v���S���� 9�6y&���i�G��"�GM���O�>W2a<%S1t�ݢ#�F�L�p��"<������z��W�^���D�������R��M����m�����W�K%U?���\'7�����I{��z���r�w�w�b��^:�b �)8���@7���<�+�D��>�oO�>��b�R�q��TJoik�z�@�=*�;��Y���ˡ���b�^���w׈�tA��D0C���l%��t82r����H"�؁�jM��$<�n�*����X����=~��J�c	�o#f���:J�YV����m�%k�!��#��%��BJ�� (<X
��,n�۝��XҎGv^⭿$0w�?g�������n�G�b������O��/�5����t��|�J.�.G+�Mqy*,d 2�|�5ۇ?��^FEC7�	��V��c"�3p�]l�������W��z�`\�z�n�.�a(q�<t�����-���O���N�IG���zH�����;O�}������b7+NQ0�ތ^�iK��ॱ
2/I��1���Xe���g��c@���8�r#�t�>C����hp�UQ'j-�o����eE�,]����]k����iѕ	�ڽt=�@B��6����I�������_��tu�_C�i7����FJ�o�_��A].
�[�cn�~�Ro{a��f´�GNӑ\9�2��]���p6L��3��+#�~�+�t��4_@9{6)�)}�{�zO�d{/1�X�A.0٣�0�l&�H����R�Z0�K��t��&$��SU�d敜R��F�lﲤ)<?���N�| 
t�ܱg�i�C�Lx���zˈ�K�Q�e�q7�j�C�C��"}G�`]���l��F�^�H^{T9j�l�������j�[<��{/=����O���j��	��p�QJ�*�G��DT��&�/U���6�8�_/	��l�	���_�@��*�����B�1�!�^�	2/�wLq7n�AN�4J�;ӎ�Zۗ� Z��a��~����Z[I���#��kmk�М��L�j���^����S=�Q��jY�R���qCK�BK9��IL��}>/�V�1��{�SyE& �s���~�*��]%�a!��q�-��f-�0�Ro�SW��G�P�R�A���e��y��G�Z��Ŝ�<���d��Jl�M���}:Z���
��@���3g�%�q�	Pʎ:S�<��s�Ҕ���q�hNOwne�)5��a��tPp)�D��ܲ������K���	�쳢A%�E^��O��;ek���9�����Nx��C��b�@�L���I��km�����s�����@�Dl7�TA�W�y��^ � +L���x�U!2�6�Y.U���ߜ�������Ao��-�9�ŝ e��i����ς� ސ��l�<�%� ���#�6��o+i@}�P�a�կ(Ro{����-�
ua�[��@BC����k~tj�q<���Z�4@
x�y_ ٻ &|���ɼ.��-K@�W������cR�%��*,s����(�`�8"�/\>h`@ ���Ȭ���Y�s'g˗�2��6�c�c�I.R���&�0{g���R-<u�a�kC�Sޟ{���	PT�nuj��p�f�u~u(�	]﹠��T	m��%��c�������49���T�M(g#'ޗ^J�v܊:����j
 D�wY�9¥�Lr�`�4D���&�{�JY�����P�5�'t���x�0�.�0ʑz�;��>^)�PF�2����^��b����ঊ@󫪦�yO��^t�������0Q�+fU��B<�?�?.SO�x-�_	`��IMǌ_��L����B�齛`�~�I�<`�d-�)i5Rf��0�����4�,U┐���#v���	�N��u������T�H^��O3�v_8�A�����Z7�bs�����^�0B����Ӎ�����-��m�%��T^!�?|�
�>Z4�����U-�k��	�j�7
�(��K��F�|G�a�J�[Y�w��X
��\U�"�ކ~���a�9��n�~B�,�QdO�ø�2����d�q�.3�ӷ�7��/����y�N��L�8.W�%�i�K��|@�M6r�	�g�ǻ�;�%��������"5w)�xw�uZ���Z���w�ws~�J�����Y�C���
���f�bn���b��^V��_��iBK<�� �A6���l2p���,f��F$��������cU!E�Gq��ݳ�	������b'� q@(��rK��@�ж5'��}�̨�����>s�a�:���ah�m-S9�TNvb�&�I�w5�a��P	 5'��ђ���R�/aoˆ�fM�< ���.�j+��V�g2���`��Q�̄�/�lS��]�[?�*D�s�@�owm23o�:0�q�!��,k^2ZM��U�X�W�P,;��]�H�_~�c���LE,v9�Y�٥�ƒ�5/���K������p�c�)t�hhTܠ{�1�Z���S3|i|^5Mtۜj���Ǚ3,6�e݄�!���Ԕ~�Bj�9��eGA��ؽ��`���co�)�\;V���El�괄���D���rdF�|_ԕ�0�&�:�����t��c3�m���H��%\��3�ߪ�x�����i���Gx\nv���u@՟�h����(*~�d?���H��'Tw5�|VQm���$.��	�K��h�⳱�例��[�ڕe��,�O@�8zD�sg.o�J>�'�^q�9��0'#y:�3���w��CuOO`cg�|Fs>u�$T�WF��	�H����E�ƕ�[����cZ�vb��c�M���"@�цk�N�M��D�x�� �	qu|Z�������=���%�[Y82����U��]���G.��SjFl�6�m�@�Q�L6P���ta.RA���"�^?8�_�����k~B��:1����76|V5����)ѱ�� �+*E��HITv���$d�3���L�oP/ �X� נz�a8ȃ7x��o���a��A��[���tc������ZF��M;�sRs�u¥��|�?M��#˴f��O������i���y�x������
_��~;Bڄ"U���z�M��=���� s���Z��\�#lU����5��"�r<L�_?H�0�?Eu�#��X�]�SHϬ�xHG�roj��h6�4 �AnPn�"�������_�"�]AYTI;!�X���n����Foo�fA�$$�aҪ�	xD��������Q������~,C�Æb�@��J�+�?7�Qe�R�"�^��F4�B'�qx��Bs����Ⱥ�z}��5텡�͵��<�M��?�L_�}��*��� �kf*�r��Gu�4��%��(�0����'�摗����O�+�r�,.S^5��;n�]�h�Pi�#$V�0ks�_��(Ӽ�w��������H!�L$���;�����UIKZv`Y3��-Jc�Jp�����}ˀ ��up*(�3w���G8��/��}�>K���}���a�� �|�<H+e*�nPpȞs�ڈx�8�D����L�g
܉5�����jn����V��-������r��#�v�؁)༮���0T*���F��pJE:`�DM=�uѝ�����g]=TÍ�P��ځy���_�܋Ⱥ&Z
���DQ
`!��8���C;��*�;.A(���s��8��A9���emo�f0F��(/��C�����F1Y�.���WBG�s$���&��X�u��p�'��X�݂n�<�8�l����d�o����IBu�/-�������	m�1H�	�i{~J����ҭF��O��,_����0�1�����Ut�NA���I��κH|�縟*�R��X��q�98}�����qj������1�P�N��W���.h�S��P__T�e�|V���!�I�B��E��}�z.'�U�¢D��,=��J.��c��|a]��/>x�X�F��=O�	��k�Ù���M	Յ�=��V%,:%�wt�˱I.�Um=Q���";�W��5[�6�|v	�[u Ow���z�|�YFO�{j�΁�#=V6<�2-,�[�1���o��>��3{BQx%��0=L�&�-h��������ע���g�ZƵ�XE����숴��!E��t�}�����/O�1��}�d�P�S<�L��qC�J�k��׵�P���vă��S��d�B���G�=���^7�0WGM�N�,��o�z����N���0��+�"`Ƴ��� ZU;�5t+h1 dK���¸�st�w\����҅�Wa�ڝ��Y����hV��o����^�:2�&8x��H�m#!�Kx���!��#�����ϩ�_@2��lf��~ �>d~p����7�o2KZH >��Q���By���h��jӷ��ھ�h����젬���S�1MV,��y��[sQ��a�|��̛��j�A@W���t6�q,�t�U��EG~��ԫ����)�:��*I�V�yCr؍���V츄v�'i0/h��S��#(�u�%�סLXQ��� ��
D>%�}���L�t�^Q��!Ͳ�������-a!�ܖ��3��l�r�QcX!�}y[1���q	���H�d9p��#9���4�����x=i [�N�T��ش�+��L�W��sF7*��]�Ӕ �Տ ��o�[˸i�k��g쬚�@�k)�Ӭ6�B�R��%G0�qW c��f�������&�+0�,+�(TҰ���g{�mߺq�T�g�I<��q��p-T�/�bԪ�?��H�7�d�e��5=�(��� u�!々�cQ>CGL����oeizt%@�F�~�ޣ�~�M�:�j�2��Rq~B�����7M>:��D��iS�L�����UN��>�e'h*�q8V����}b~��nAF�bB\t	�'�g����G�sX�Ks��;�W�I!waJ�j����� jύ�}�e*a�|�k�a��� ��`��tq͈^';,E���8p�&��"8�~9׌:�Aa���:L|g�5O���E�y��S��ޞ
5s4�R^����@˚���sa�FWwqz
�8U_�
!�6ur�[3�ɱ�%�ji�)ѰBZ'�Do�V}���mGGop��������d�- 
6����s��u�m�L��Ы�ZD�w˸���~o�[���f���C	C�����M���&'DY ��l5�"�?c�Ǻ)�~�K��2Fh�h�g��=+i ��3��´��[��[J~�����+8ɬBf;�����:�S+�U�\4��'XgT)���ڶW��Fo�W֕oB[�����]��3�����JU����\aiΔ$C�)��]�yɷ&%�e��r�}��B
-�|Y*(@��(3O�P�%�Q��_S�?m2�K��LL�(�I��&iµ��Q���e���}&=
�i�.$w��8Xt	a��c��2x&I�SRM1�6�0�rM�4�J��`EUF�Y��p�K�?���^]���� b RS$�ܙ��J��_yaE+�37w��I��*�s�
������QDi�R3L���]9��NJ�G�-��`�s�-T�~ �N#�582�1_�֏v(}f�^��YZS�𭗬u{N�w/����S�l��ɇf� �u�-S?�rB�f��¿,����=u����1�^>��{pٝ�ͧ/�ܔǈ���^T���`��_jr� �=�Ji�I�ܿ���iaҎ��z3�-�2�<�n�G�0L#�ф�S&87䡗�Q�2�M�P�V�
$e�k'�}G��h�&\>�<	������-����=�3#�7������U�D8=�@tr���]��ϴK�1Q�?~�#�m�$$uj>Ҳ���5�ƶ/��(<ŧ����4��*�!&x���|�[
�50�@U9:�1�)]�� T+W��>��/�6��W���k�]���z�Ul�f��p֑[M׼��8缷�P"�$E��?�ǽ�9�s��_8�e7����e7s,b����	P�At$%�NV�U
n��.��H��Q�a�4�>+���#6��%��.E!w���O$}��E���#��G벰3�����D�]r&,dw�8Gެ�Ô�I���K�o�T=��|����6h_ �`^i ��|�7�O��D��cS��G��E��*���,��x�����t��4���;`dV$�b��H��8"���Oa#'�h����N���P0Jou�,W݁Ŭvhp(�G͔�@�kB��D�5���K�BAh&^��c6��9��`� +�3������O�]r�81r��1�y�i-v��3.-ڤ4�����n=d,�L"�ނ�o���;���S�~��\gW��NWK�.&<��r�m>UF��&.Ӡu�mt�����X�¤1ɼm���Y�f+|��"{X���D�B9�!U\B>�am�W�Kܢ�ᙠ���Q��]ć����r�����}�-߀�x��ຐ�^n��~�A�z�
��m0N*�bx��u�z���W��IBr�d���!C1j��Q�����J��Q��{0��=���O��\�Y�w��7�jAEV�����N%�H~s9[C�qT�u�ą��4�����д�ߜY�|Jp>�s�4�E�Ldu!�} ]�C_�o�O!#�&`�.������l�R� ��`U"Uo򩕊g���#����_EK�Q#���9�or�G�lU'Q��??�j<N7:Ό4�!X!�.v]���g�W8�z��z�x|�!-@Ǿ����#�xk���׾���s~�=�ڌ	Wͦ�qtz�0@n�D���|ь��3����B�87-�t@+ڑ@�j�̛S�Y���b4�����?�h��n�)��ѣN1:e�E�^Z�y�	��X�!1��y��?xh��6"��JՏ��7�� TH�(���V�((O��|�_�>�ʨ� e��k�o<M{+Q�?N���I���5�p�����Nַ�0�[VSL�eO�}�.K��0�BY+Wٺ�~���P�g*�Q)	ϡ��Lar7'��F ��=M���$�H�� �/w�e,0K���h~0Gd�V���hq�iDl�-��im��hj��� jp�v���SJ���X�x��N�Ma��e�`	�*~ǤC�'����ˆT8�|���m� dʣ��-�o�����'��vM���۬Є�Pu�����:�>��j��!���ve��Kx��z�Nm�Q�ǯ�������.�1Xl:�~X��\�_��Ս���.C5�^�,j��+R�2h��Y� њZ_w��PͿ�\��H�����G��,�0�K��%�/������B�w~�<�+���TzL�������-�kc�<��F�SZ��`KnM^�P|͞��������Y���T�D��&�!��v��4l18n�#�-^	{�5�4�DvVG(I�٦�/�3j<*;�NEL�GZ#��T?(�~�r0���:G��>�Lg�@�Ny>!P7�=�ƺ�JV���o7�Uf��]\��N�Y�j���RG�,a��]j���R���%'0QA�n��&4v�?�o�l�=�/�?qÞ��i܁BI����VK^�fk_V�����7������I��������Mz�����.����9�@+s��Y�p�� �V�ٙ��q�0>�3�}�'�%�"�/C@��"K
�|2����	*P�����W���%o�$�`�5G9�����8#���#�/��#*�c�lVF��<�:n��Au��z����u#9��3�)^��0D���*�K������
jk�y`��⚉o�>����r�7�;�S}�<0�j��wE����0�1�����%�aCkL�`�0�9'��m{?�5�/OB��0�_��_�eg���i�'%tv��5f���>)P�L�Af؉xGz�J�5m�����<j���{��˝�j7�l��PBB�S_�$���<�LP^aN'˨�3�z��iL��õ��������k4�7�-�E��z�"u��\��_�A$b�>�Ʃ̼{1ބɉ�J�=�L�֣}c���\8�#Ov[I�=��b��%��Ktى��&e�_'�W�K;���i��l�
q<,У�|�(Phx�)�pm��%�ѻO�uΞ��w��o5����8W�RB��~2�%uM��	%��}w=�I�29��;�tQ$�E���~^�����a�IY�{�Ѧ�Ī�m�oJ.Ǩ��R5�3.ۏx y�n�`����.��xZ�W�Eu!���2��O���}p'օ�]��g;S�h�JčW�%Q�+9�BO�-�;StI���fw�Ċs^=(H�A��r%�o4sW��X76��Y���uG�Q!�Q�ԭ���S
�5��x�l�v��ýܶ`2�������+78�c@^�1����1�fG���@��I@S���s�����@!�ھ%b��Ɛe9w�hLU|�_���]�4K���_V�-!�q�P���`?�R��%Ϥ�����%�A�|�P"���J��C�[���O�O��XQ����Nd~��q&C`�r�=��c��M�$��ƿC��)Ł�u�Q x�R��;,=�kvF06�M�YF�Z�a�s�0�c�Ȟ��IM�b��MlaHv��f����c4�5Q"o���B͖g��kдA��"�_	�X��2RGS�sd�H������8|�nj��Q�K�:ZO!*Vd���R���S��5�5��h)�4�?���Z۵�OaV��#���衑��VC�X,~�.^��&����ά�	��ݻ�:�#�b�bM��<t�྘-o���4o��4�C6�	��Ƭ{Zg��yg��ÊkjS:�d&�K�_~k�հt�6�d��:JcKv���|>g)������vm���5n7>�U�ҡ7�PE�@�gjS*�������
��R����(�Ň�H䙘^�ϩ.
�L��Q���&��Z(U3�r��w�X`�
�c5�׮�+`f�)��!@��[��˱sr��m�,x�9��h�7�c���e�6��9�$��?WX��|�s���[�d���_{gL�!���5���Bcs'/��b��YK~��#�R��&$��Or�ENt������s��wa���,�A���*�x�`,��l�T�0���~���d��W�]�ύjnR8��WU$��WACGO�%D�
Bl�*��e���]�聥�Z�is!��c!Z��e���.���ݎ'��ԗ^�.��'E8�AG�
��p��H�W(U��XO٦$��f]~��3��B;��\��g9�K�nG�\>,�*'[iA�H�(�*��*���q�ѦS�ۂ��.�l\#7	���G�W�<�N�H�A�<�O��M>_�oN��4f𼐭~�	ү�n]&
�H����L���Ȍ�ϴ�����1���RNX���G���Q�ƻ��~n�ai�*ܠ��W
ʸ��F���D����C?��*�3�#��!�t�4t�y~�(�:!�Aw4rm�x�)�֟!� 
jͯ~nA!i���&�/s�+���Xy�5��ޏ-bЈv�u���;3rxmG�Uu����t����BE��d�� �����=p�d>k����X���z�C�'�����Dv��5���mm��'+9�-��_�&Jy�ɜ�,�;���!�@(��y��it��h���=t���Sh�=�Z����폴�ʶ���+k��:�4O����s��3���6k������<�����o�#=5]�ާ�4�Q�-q�-�_��QGn/#tk��KM�Q4���s|fOw�[����ZpN�q��AP<�c_/�ҷ�=o�&�`�]	��������lm��0�,	ƻ��a�Hq��ׄ�Ko�߅|����D6s�(,S�a^l�+��?��oװ^4)�����QGZj���Ù�����Մ8pn^� 6zL �5W��6q��j"y�F���2oȱ�&k����As&S',_���)�6�>�ڄ�l�yD���#�&�\�!h�����G�ш��Y��@Si̊��k%yIϜrPB��s�A}1��Z�Tn�E�y�Ü���utBS�`��=�pZCQ��mF�F�<��*y��RhS��w/��*(;o����s�bJ�'G8e��%���G��.�K��K��E�4��?r�LP*=��5�/dͪ�_^�
�׏����8?w%[�D!�0�-��dV�'"�(^�euO)�0�E��yk1hx�=��FＸ-
ۥ��X��Fqb���	QS�`L=��i��8��~�@���)���t��b�:�-�����2��
�O�8����s��;�S�,�[�ߜӿ�h�M��Q�~$H�u��ٗ��]���x����;�'�޷�b�˳ո�L!!:*c�m��O��<�҇ĕ��]y"�o�����}j���Wb�ɺ�%���<���� +p����i�0GSx��"<�>����S���~�N�p���)�V�q��ت�!>M ���}�O��Z���*�&�
�����1��E��;R+�8D=����$]^��.Brذg��@�΅����|��Y� �%��B�z�C�
rU#���3+b(�,�c�8�c̮���k�T3ׅ��َ������9��65@���P�>�XZ��'u��M�?����ǝD��Jit�N�(�i���\"1���@�A}ۋ��f�|.�y6؎ǜh�z�>΍��OpU��l�f��R���e�ˬC���w��Mޗ�C=B�1dʓJ�h ��vF�q!����)9�Ŕs�	3(�5/�,��L:qA���
��.�� ������t��#I:2�uvG��40j�$]N�Τ"�g"���Br����nN'b�#e�w�r���˫H��E$ë40V���\�6���;
.]1�<"xژ���dwԹ��f�j�Y0}<F�Z�}7W��smԫ͹D��@���7��Kt��	W׌_����2�ʓޕ��P�0Hd��\���+T�$sՌO��N|n7Y����kP�Op�Y1���0����2`�g����'R���A?Z,9eh��~�j#u�^��:6LF�����ģ��M���� Y5�|@�9"��-�;|�Le��\�Df�w��}MS�>�Pa����!�A��b��~s��Anzk��@<�$�6M]���k$%Ԉ2�a�/ގ��z<�͸X�Ԏ��Ж]B&n^�S����ao?L=�k�����0�~�����COtx�f�Ԍ�\��gK�Tӓ�f؉ں�մky3*�T��=�.k�B�۝����?��dәt�LP�*�-	h��V}��|ڎśc4/-����f8I�ć��S���e��v]]�L�'�k�r@����,_��1�W��I.�[C$�yG����M�gVԙ��doS���"�a[�	K�Bt���@���|8�l�)�*T�:�$������g%�ZaD�������-��"�X�%;����]`&���l�!Ձ�V�xuK	�tt�,Q���֑dn�	��:��<���q���l��C�[U�p��Zxܿ¤���������-����$��i�,�@����Xu�{������0��_���*r�ų�p�`�p�W>K�P�cqQ��N�����.:TP���s��_�f=�86J�{��my��`x�mQ)���f!������"b��C<-O��W��n�d��*�����*쨵��K�J�6j�DT�.{%3��m�m�KПKB��(o�-�y	�p�~��Փ�c�<IA;�2�@L�������s�,V�-]�PϳcAEa��<m_�sk�r�@�.NS����p��F��L+1ί���x���?T�a09PRb�q)l��?�u9��C�/���A�	�;�l0��b�)_!�6�RZF�	�,�����Ù��E�R\~�j���{=�L��P����R4kLђZ{t��=�#]��ɰ�~WYw��_�rZe!�'iM�G��5�n|�g��{��"�Nx����Aic˚�h_��H��U�<';a����$t��<Mdt^3'����\���ە��?%]��!��q��/�m�a��t3U�i��E��Dryw�mPi��I��|�#v����Ao��A]�@q5���'@�v[!G���t#�=�,n��~E�����|tBdt0� ؆�g>x��Ԭ����TgBRG��R�2�����?��;{ef�WS����'�$��
�E�KKU��7͑�4Y�}��	.f�[���.���!gq�������>�d��'O�JN)	�#4��g���W�L�4c=����j�����/Δ]���Y��(��%&��pd��R��J@?*�a_����u<�2Lױ��8�3��χC��TV\+�3`����I���d�`��J�+3���Z�t�Vu!�~Y=��� 4��Fv��K���4�l��\5=���*i�w���[&]B֚{A�5=G�<m�!AX~;7��*o�w�gB��<�ZY��N3|[�k������Q7��$=�گ0�z/��ݬ_���}�ж	t���f�ȟ���R�J�3�E��ۢ�T�.˟���At�%�v%��0YY2���B�&�h�m�0uX��0\hu*��2��Ƹ��[v����m����.���1/q>Ӂ����_�_Pu�"��4LIa��@��Ȭ �}yIqß��bJ�X�0��,o�����3����U�.���Nj��>�����|�QE:J�KC�k	��&5�S��	�ǜQ��э�;�̕M��,u^��8�1�R�\��p�4¼�t�$R��R'��{���e�꛳�N~J��O����q���#�r��	W����Xt�:U���.A���=�B����NXY�k�	��o	�El�Y������9��V�������,1f4
];e�^�M�Hʥ�M�r�Mo�l���uCa�N��'c=0 &��5�di}�#�����f���:߫����	�F��b1��=Pg�-�+����T&l���L������7�66����j)�y��i385��]���&�@�i-����5�пQv�@(��-܀o���W�#tE6�s =��Y'<��̹����0L�<%�HO�JZ�G7f�r�gV�xz�cR�ӶU�h�\��6 ��PȂE���X[tT��v�'�܄ݖ2AY�5{�M�^\y�s����*�E�o����q�Z,�����\|F<����GJ��;��K!��h��X�e�)!�n��"Й?!1�������Q������,�2;@Mʳ �(J�?t�HO�t��|,�U;]'ޙ�F�D�w/#{Ez�v�?b[-��ۥ�;��\��W#���,.���H���X��g�W����}���[��#��f��o�!�./e��}6Ɲjl�)�7��v�l����!�w9�����O��R��l
�|��-��\#�
��_)��A{\��w��,�~�_��RSp��(g�>Uc*LN3�ХWZ��x���O�G�!c��@�����|��W�t��D�U��4[�
JY"�\�-Pk-�C��ќ���;U%�/��f��䧻3tB�H�1�m�*ݣ��j-�.�U �$&�s�45��[�n�[^���N�A���|/c��BR=�.iDU`��B����(��^�Ys }Y��2�DP`����c@N�a�k��,G���?�����H���-o��S0��33��{�����2kSO���Z" ��GO�ֺtd�\�3�Yi��&���	LMJ��ѹ�9FW|Ll�i�n?��Y�)Z�[MZ�������S�߀����D8����u�6D�����W�馜D*L<Wq?��g��)��]��\~tcǎ����ٮm��Μ�]+���W|���ʴ%U�H�Lz�F~;%W�).�@�������k��12��8ݻ�b��ݛTګ�٭:��2P��/�@�6�$�}h�$�p�����oy�R�,���c��d4̞���6���Ë��ָT�$�W��p��8���Q�Ļ�"����P�}G/��e(.�K��%( :rrhL��ҽ%�ǋ��8կB�*َ�Hy�E5�+*�FJy=����(�7i�����W��pj��O���$`�:�g�Ã�^�6}���� �b?ve�38j3*�����&��mc�I�+�04��}t9/�������O�;��*�;�h@8�>n`�Ά ��0Д/�������N[�1x�$�ad��R{m���D����[�C�o�@�ܸ�e��ʸ���4۱�.z@�����.�^��a�i� �0kJ�9�nM���'ࠡ�<c����$ЈPU1�[�ޗ��NKw�0�7}J�?6���2g
�=�(��T�4Dΐ�M�aN��Y��K�3.��D�I���f�n�����3%vYK��ʢ���C�S�u��!َF}��@x�`��vL
K�5�:�8�����3��
:�Η	�T}�N�����z8����ڳ����n;���\��i$�ľ�BB�h6D�Iީ��s�wGJ�ܾ�բ���� �<���n���R2AP�r�Q��������5&�!M��m$W����1�c߆�\9au��z�ɩ��몪���:�ȓza9�����e�'H��W���'Sf^��U��r�S�"��[�`8���!>�{$�F�Ee��L̉v�T����,�-�M���s#��"�I��-3��0����o�($�0*��o�2Un��T��$�ߍc�YhT	�&�9��v�Y����Q�	'��f���i��X}Xm�W��)�l���S�"BqjY
�ڕS�JYc��#�4ܥ�'ܗ/��/�y D�t��Ŀ�x���������0��� ��e���F��l_��Q�H�$Q$�>��L��2��L�V8�%��B�^����T��H�G
���w���k<[��j�e���m�������W�r����c3����9Մ��O�� ��e9�x����}㢘��]]�/��t<����%����q_�ԗ!��H�`�FohGu��"�	y�^d��+�{9k���h�I��ƨ� C��U{>:����-�����@H�� ��_���pݾ���e�����#<��D$�����>Ts���`J<X^8�oDoa�$��Z�S�V�]I�L�F`�d�7Y����gy$@���03@��~�8�Db�T�j�����Ϯ9��-�_�����JMT�W%�V�Gyu\Qm�>J�f�Rm����A�:I�����*��v��څ�\���lJP-��=��c/v;�Xm
��`���ɯH#�Tf<��s��T&c�		�%���c�z��Š%=��U�����M.xC��ǻ?�.r�5VX:P0�7v�`��\��_S�e���g�	?��Ʉ'b $�9Lqj�Bk.�1��*I,	���A�z�<Խ#�Z��+K�U��3.�5��c.���=~�d�D?��<;��W���	 ��o3���!�ՄK�>8�Ĩ���%ExxR�PC)��p��F߭��I_<�؇n������q���-Қ�t���3{ʖv�5d.Y�sE��n���bz�L���F#��q�f�G�o"���j#|
�w��k�s���Xa�0M�zsP���@�=�:2���x���EѱR[���lB���I��0P�m��_|�<���J�jE"l[�WF,>��L�d(�F�B���1\7��@�	�gjD{�n߽@��/��҂�s�:&[���t�u\N}�Z u6�^&6J��)R�gW(տ��!�]��)S�:��۞�*s���]�P�ML!����0�'�3O���_'J�Gw��`D��V��[$Dd`������X�D[��K��y���jf0\�B=�XC�`��l)�����_�����ZR���;A���k`2���E�&��xp3�,��h�I�=��^^��"/��L2	p�վN�Ră;Ս3|�w9�۬��C�I¹�(�!ۨJ��D��+�����jz)�L,
� ��Ԑ7�>�ɒwp�#V=xTP�V�w�Ia�b�ɞZDq :h��������8��b��pw���y���B(	�K4� b�� �b"�8�V/�23��5���U)��++T�J��]���M.�רц�C�eȸUU,� Q?�.bh�7��o���	Ϣ~�m �:�#̬�Y��?�쒌u��CP�hΆъ��E`�R�|S,���tI�v�sc�h��B�6"Q��-֯�NjW�ϨY��a����L�܋	�9  V|K
$���vT�B��\��� [N�E��zrU�0�ʆ(?�_]��Vح�a�G)b*�8�i1P�p�#��MC/o��MF���V��^��;봲F��B�L��7B�Ƞ�d7C�����Tt�63���e؉3�|0Y������%�0*��ӗd�2�D4ZA���'׸&ա���ȭU0�؝8�B2�7����̅n�\0�\?�:�6;���N9�H��{�PG%�Ք�w��-�&Nk�g��Zu��U�	����`���DĲ7�%�B�N�ﻜ:`�����5D�f���D�!Y�nT_�겚�B�"�?x$�����H���<�=O��\�wj�A�L���`��j d��W<Z��.�E��瘩��55!�u'g�u�P'���	m.�v��汛zo�d7��JxQ��u��%J���S���_�O6�A7s��͕7�&b�}��(&�'m�-�I�������/"nb�Z�I�"��_e�'�w�j�� ��6O�нhSC��H������M���X6l.<�rd��Hˮ��
�/F'FYq���N��D�����Q����	�/@g��<��cљٵ0��mu�Y+��R��;Od6�T�F�6���k%ה������,TS-5+�<���r�
�U+�֧�b}�?�~��V���T��������#�K�c�r����o�#e-7��%�U�~Ĳ�o���,5QUFm�=��%ڐ=�X-v��FS�X�;�e��@S�$e��&T=_w46"��hh2S�&{Yb��Z��%�$d�O�Uq�P�UgU�g���ZzR�<3�/��E{�&�R���{W��V$� ��d%+�Sn����h����q��B�@iF��^��yR=G|��;D!vm7�
�s�|�|�^>3�[=�C�E�=�M �� s w�����b_�,ʹ��r6�@�j"%�ra)�1)�ia�Ւv�nS.�,�
���ѯl6��b?��}�<��"��[h^a�%��ɀ䢇���g�W� fԻa��T�D � �,��A6�G������?��#����j�Xr xz�.�{�@��^E���9��tuˏ�o�$S�~����٢�s�
��a)5�'-�d~��s��0i�sV'��v.t�VU5��Š ��#z&��b��07%F�O�YĮ��2S�$D�/y,s�� ���Mg����%	�OQ�V�<
�2\�`-���~��cz��kVS�`�=菀P3!T�%�F�lk 8����)���c��!L_Rd�#�ŅOs}�%��Z���6�]�Fe�Bdz��,�E� ������A`w�&i�����է�_�yp��}�(کD��Y�і�"����u��c�zb��+S]z���ЋW��kh��a�m&�n��%hB��0ˠ��y��V�2�"Eb�'E����-�;��.�r�o�r2M!��*�����-|!��f�ȁ��9�K�܉v���c7���Djo]�[��@��3SH_��U�
GG�>ٮ�"/] ��F�tB?~�\6���0C&k�����ipc��k�����A��d<2���˂�%f�0-� ��U7LF�N�
����N`�A����S�}~W!L���&,^}���k�S�g!m�sZ^*Z�����9�]�##�Og��Z@�@�%>)(�u҆Ǫ�\Ox5o�x�00�Ŕ�a2����최p���
%���1,��o�+�b��!����:��L��8�6��?>F1օ��x�t9�%,Ӄ�OW�o��3�&RYy.EI����h�Q���Ct�����9m%���TvV8@�#vv���W���ǪE�3Ը�yѰlu��u��Yh�^K����>��M"��C5�I���M�5��f�Q��M�'�O<�eޫ�z���Ǚ�|X���U��g�)M&o�b�����/��#˕4�/�O�t"���\CI���k�A2��c�~��]6sXl�z���=�ʰ�22X������w����)z��Rg�G!��nj/��
��o˿��Q���:�p���ʍ�(Z-����s��h~eZ�2�w�ڠͧiGz��VW�#@8f��wD�_�B�bL8j&V�s���Vmh|�᫡sU!i�[=I./ �'�MՈ�&��Ӛ�p��@��#ֽB�;U�z��I[�h5F���'���f#�Ŧ��)�S���.���l��Ѷ9�e�c�?�?�ߘ.�J~?@럔�_��"�1���+��%2@}�x����c�Y.��)0���VmG���φc8m�Iǂ��`�մ�~2��g��Ԝ@�7.�DX_�J܍u;�-��;�E1� �|�ii���	E�E��6J�<�|�kg#�q�C`'g`���<��9�`6e0��~wqM� �00��k�4Q�W5�,-�}[���j�{6�pU��A�&�?S~g�#��~+oo��bM1�<:�������:AѸ2����7���[s7�]��*��y�tx�,�(o%jd9&��o���QR�0U��+�l�GO������rQ/"~��L�|ڃ�;�XՍ��,�%� �o�w����lBq��4#?��9З�WEM�)Im�e����b�bj��m�tѦ]j�#ۋ��\H1�L1�HI�@m��"�#��#ʑ�pP�t\m�V�W
�լW�����v�wݭ)�GB*LR�n4��_}��r��L���N�s]�!�+����ABz�7D"�m0[����EP�*�oR&�'�Bn�X5^�Si!d�GV�F��;��*��:c��ݹN�A�q�N(^�px$�i��~_�D���\���������x�`D/�lrL1�\دI)���y��ـ?��:�Z��̤|z�n5tl�G�1D����N��ۢ}GJ��j�h�ۏ�	��i�=1�;XX�,��G��iaز�� B���[��d��bBRi�>ߝ�n)��V�V풿HE��ȼd$����FK��7���f'�G]l�==9szw��8�[A���xup�?����|2��~*���y2�z�&�e�,��׋U�hy�)hڌ*"�]�I�����+��Kv�� �l4iPy��=5�
��/�-qģ��;�}��Z\R:^�Mw�J���^���x5�;��*��֎.XmNH�[��$b�����o�2p�[q����,�t��ctl��9��]E������)���Y��qU��9�r�s�I.���X���v��6���e�u�����R����Κ��ʐٵc͵�H �kdt*)ă2�Ƀ}��ze��#�Ix����"Gk� �I7+/.��k�$�G^�O���,�O�(��c��;'��޶�E�(�ӻ_%�M��!��~�E1%�{;�!�dN���I�O�{��'X�f��]��o�ǳ�(ג+�wǱ�PLȃ�+I��砹�*��d�������o����.<�:��õs���\�m����Q�\|V��b��jg���� K���{Bʄ��~�d�Z��%�T�^�E���:����|���]]U��&���-��~���Yz�����qձkd�3u�0v�,��v�pL�R+����!^��*�R{&{S���ێl\b�0LM�'<����'��~�g�hա�L{�����N�؍�j�pժ �>�fJ��-�"�&f���Kz�Rx�X�7�o���R�;d-�{T�/PR�գ���3�EH�7�m��9�6�U�m��>�<�� �����c�A��K���p[����S���}�3BS�yݝ��k����Ha�-A7Y��ji3��t�w����f����A:|tӄM�lL�Ҝ��A���nQ+�<�/�[t�}ߖ j�}�NJ���#Y�4ɼ�F�w�(6�.)�Ok��fv��-�_�	e��h�J�3���r����,��(��a#s_��7����|>@���| ��$o�,�FM�ς@�C_9�|W�8=Hة"	,�ث���}��ї,��*�М�/��ɴȟ�AQ7�2�	E�{f���AX�|�[�JɃu�{�(\�|�4ϐRf0�^���'����4-�Yb�����- I�!f2&>A��A���+� ��VP�	�X��Y�v�k[�;a�2}U�v��Yr��s۳��m�8�3a�C�Ŝ��ݽ�{�&$�i:��weS\e�0�up�٥�܆N�r��:���P?u�)ZM⿃�ۯ���Jg��]��^���k��im/b�x��	���Mf1>z� �#mL��C>U��T�H4�Hs4����{J�9Q�cts�*������P�ټ��!0IOiU�Ez~E�$u���8}sp�y �Ekq���#D?��c���
���I�H�_痎E6��4S�V���Y� Xp쁋���419���KS���0TZ���W��I+�i���U$Z��K���槭:O|�Ȳ�W���g�|9���`d� ��ƐKF��odn����~�҄pG�k�䳯Eiy�L�����Ta��㓅���ojᰋ>5�Ua/��#a2�mMt�hۦ���Xr��Iɩ�zX�F��
?�{/,� �N����Ņ^&"\tI��|�ɂMn滾u��-���{|$���Zj��ЧP��-J�{�!��0U��;V�_i<=fA���Ɩ��(����,d�)���W�?���RF��-��H��삦G�Ww��l=���5�y�,��M499�`}�G����G�y�_���&��a�~��������]T��!��iE`�p5a#ո"I{VI��G|+�6��{�0~T�i���E�'VL�,�X5�14}ˈ��m6 daZ!�O��]]���Y���'�"�%k�j&�0��H�y��Q�i|��1=��a,���,�QR9��0,� �i���? 1vx��n�\�ߌ����.e�瘵s�2EГ��/<��_����˭^zu�<vKh<6����J����˚�TP�Iaԑ�łL5�kC���J���"�2�h���X%����8+[����.���7��\-�og���n��*�D.�(_� �0RQ�����?���3����IʳG�cQ4<���i?����M�N��r˧%x�8c����nngP�g��Vᛧ�0~ۋ�}�d6�o���R��-m������dĥ�#�0k*��R��Z�V:L���bJ$���_�Aا��� C�|���,w��u�Xj���w��F��hi�<I��-Q4�k��l�����C xl:�$�<'>��@q�1F�.���p�� ���(&���=���񚉨+�Hp~Ƙp����t���LA�9V�����~�>Zv��^10kb�ꢀw� �[#��&;��-�&H�81"OP;���iN�n��J�	�\l�R>�ܹ���"*��[l���[���L���J����EOL��q�O)r�N�ui�0�hH�����o�{	�k�����lF_�g������pϛs��fֆ�&��*�f�>�ɄXI$;Y��<-+��I�Z�9�Q�[A���[�]��,�w�l��!+פ���i��<?{R��!,ߒPa��F��ϸ���(d��к��Cp7�>�����P��o���>(�QW����ɦh�[~�1��k�V`������o�o������T�Gs�J�JW�$Br���A�t�YJ�X��I���
g��R
�t��o�'�5AmlyH�ZW�U�c��Ip�c=��V5"j@���?2e�A/�h$�$�}����4�����)I�a���5�b������[j����"�0������tu:{Ʊ��9��L!b�)A�W>�4�rS��<�R9��1��f	p� ��-�L�о�M�|�T��?zic�!U��%��W�l]B3�m9LV1w;hah�f���N���+��*t=��Z�na8%@=��5^֖-e���o]`�D6��,� �ڛ�m=��ǌ�,��(��|�3��։��<{�6�߿d������)7)� k"z<	�9�}�oL��A�b^�z�T+W�f\u�'X,��ȏ@�{�6�rҪ�V��D���ղp�e����JjEf�����g����f ��۸wk�h�-�DS\�P~FQ�W<������KNÍ�^]��X@����<��a}�"
e��mKb��j��_{ͨ�&������E��˵p����pD��#k
xdBY�8Yw�E��A
<��Q�\C��P\��4�|.�<1tن��W�5�9�u���;����)�jET�X��9r�ǩ8Gl��<ȁx:��p.�ڈR�7�E~M>��B8�	ڥyG7b���͏��`��j\x�ԡHT�9?��	�o`�J�����������'3v^�P�a���$�z��-�F0���ޒ����?v��g�٠�ڙ����(�R������*��ޝ�=�i� ��;*|3p��y�ʵ�B6�\�5~���~�vͬ�oxe�t��0�gƈa������lǚC*�=���R��+a� '��$3���Pk���m��
�H��[8[���J8P��y:��^��Ժ�	��;�o�J}�-��Lc��u�Z�'�<����
��	>�]�-qǞ�U2V?_:��� ��/�K�3��vz�R��G ��Q�"'Mg�.�|���J�̚��?˗�	-P���hL~�t���0ܡz��dMF��4�Ǹ0�q��o�<���r_qX0���N���~�a��Q�:Bm�Ĥ��c�BA��zt�i���2�>`+�˦B��b�	K�5����MCZW�Fޫ�����e�7���B�������2���D��˷n��1�zzf��O��rR�ӗ��^����/�19�:�6���@�B��l[��b>���œ(���V�h�̱ ꊢ��`~$1�J�I��<N]�&l�_�)�!� t>�e_�|	*;��1�u`&�?�J�4`9���$�W�n�KNK����� �p��X�գ��3j�ɗ��&-���]�<�$L��E� �qv4�s1��Yc��0��u��^1���:��o��%�D)iŌ/��|���e�w��hf#�$E��MWQ��e�}��F_��t|�DaԼ}�h"=(�Gܞ_'�Sl��;9Ҙ?z�;jt8�I�G�>e�s�d�Q�I��1�l�Ln��c�6"2�D�����bۛ�9�p0�Ӑ� 7V��=�m����n�1�Ă|FD��$�g�H�}��a����}�����8P�~̯V�H� 2��pZ��f�KmE��=}�t����ġ�o����x�r�9qw��_b0�k��f�M�a�� x�T��V�d�ޖS,�4V@߰����f�?�"�.~�Ն^�#�� ���������)a18ϓ
^����혢��0��� :�5f�˩�[�'!b����-���2�z~�$��7Y���쮙Դx(�����ڤvؼ�[ot�D�
G�R��Ǒ��:�\s,A&��g��8w�Q8��_2r�,���IM�����b��Vԋ�'�J 7>�Z��`��Ną.a���#��j��MMK9)�1u���ϡ���b�e[H�$���֨5�V�.|D ����Yt4���Fߐ�9D���⨝�4��oIVX~��K�>
�}T%�!�L�� ��hrK|=��'���bj��0@�(p�Z�r�
�lH\"hwv�`V�p�[�M���x�$��z*h�G��C?ٔ=j�jj�^ڴ±H-2!�7�ûJ�Z�]��|T���/,N��~/��|��'g�`�����4kn��[�?��P�nkH�%5eD��,��\b��X�Xt���S7&+Y*�;���F��8��	�Nh+���V0�m�@j<B#�f�^4�&�i��xu x�� h��o�!�xp�@sC�����_�u<jXI����实���Ǟ��pb"��N����dt����\gZ��v����I�zL��a��6�E�ޒ���'$f�W�>s~��a�N�(p@��c�l�x�p�[H�o�B�6�R�!���PYNE���:.N9��8�
�]@<��338LæjKZ4����/ɔ�Ò���}�A�p�W�|�c5\KjE�"�Z�W{
8���:J��`�*�K�E�V6V��1��Jx�_m��q(�EK���*����7-q������l��J� n4�{�t��Ut��S�o��:i@6�!	r9�����)����܌��<��5{��"?j;�'���j����O1�?��\(U,U��'9��r�&�[�t�w�<��W~_�xk��&!z�j��t~���A��5��UgظЂ8�Θ� �k_Y��C�������&��3�� ���v.��G-OGQa�m״�jZ1f9$#�i;MZ�_n���m(�c�C�A#�_�ذ/��aC�W�J�>�(���N��򢘝I�c0OL6�#��)��V'�_��Zc&��6�����.Ȫc��l��Š!'�E���Y�7+0�&�&*%�&��u�#�Op�o`Ns�ۥ�c�CnB��9�20Ь�yC������8R�AX�wZ�.�~óN�,~d��=E�
�ph��6`�L��#6&��`yI^d~5�9[W?we��_]m7R}�*�� OG�~��Vz(��d���ן��'O�T�bA��~��+���#�tzw�3|��q��k�{�@"�.,���}�'����6��D�����j���v�~���֗��Fmڥ�+�-�ҧs,�#=��q ѝq���v�}�����f�4Ѹ3B�ReM���ۭ2r���mg�ıT=oЂrz�&$'J?��8jG�$;���:a���y������f�wX@�Qa��;Z&,���B0�x�u5�gI\;�L��`_�f�Z�ES2Ê�>�W�Ik?��`�k�1�����.�4�H��I�8�a-t�*�
��\���&��d�?{񋇰t�d�ƾ��5G�Mf��h��Ǒ�'�b�d�P�TH?�	i�yz
�4�P�P(��< �D�٧;�{���=Gy�S���L��Z"���by�1h�c[EL~{,Ek���!��;�' �<k��8d���y)�t��Y�w>��q�!��"Aȿٱ�G���2��DQ�}߉�N��Q����R�d���ƫx��c$]��$8�THӧ��l��#4�?�/L��S��G'�Օ(@�t�d��� 4�C���OL7��s̈�,�l�*��t:���/Ş:M��r��~������:�;G��P�]4Dxl�r�$�1D��P�����2�W�>�ؽ�_6���� ��5?j�o�%��/�G��z������ݟhG!+dk�1���e��P����9/�4�& 㹙����Q��T�\Hu����d|x<I��E���=N�fn5��"5L|�ٞ� ݕ��25jXK
�@z�}�������YV�:
��?�|�7��S� �)ZH��Z�Yx��(�);jap�r��H����)<����n{��;π��e�sGA�sv��u�0���$�b�_������I��TY9��-b�h���A9Nf�s�8m�h�����se��p�#Q�+��ʍ��%d�'�s�՘�V�u%��r�����!�_間hK ѡA�]��X�ރ����P�t�W7�┸�R��>�:���Q�Y4�����8����j��࿿�Ї}�fs^a59�SV�/,�3"p&��ͨ�&EԬO��7'v��G{����8 ���v:ӂ�0�S�Z���H$A��L�ɏ� w(��V��S�;�(�ƪ&v��p����)¡�����A+�S�xd���s?���K0�'u_j6F����?j�(ذR�f�- (����y�w�*qʵ ���\3��PbW'�=V]%��L�,�ʤ��Y�f} ʷ���z�i	�wC�������D2v�h9�����3�S���H��ܷ�Aw���ɡ�q)9Z�Ji`���T5��T��Ona���%4�A�Yc�&T�	�'Q�LKj��/�I }Y��q~&C�w�s:��޸j�V��s���7�����h~�a���6K9��bỎ7Aǹe|}+!��6�۱>W�NS���7s���KEE����;YV�EQU�{��.��J��w)������K5�̳
� ̲� ���u�$v��6�zӖ.���ǌ��+��kLW�<iM�ȑ��K�^��E�����x8�~���������E�?Q�A��r3�v�Ɍ��9�Mh�z�WmX��_<���fBa�eNH�,f��pjN�r��6k��9�H}�RpB�'��uf���`��]�K�G�ri��ލ6�sԣZe�y@��W*�6������o�ԕ�2�Bp���,������+�J	��V�%���-��d��U�����R�(�x#�E{f!h�X4�r�_��Lj�27$a�WdpM�S��^�ן֚����n`�NL��.�=���-�w����f�8�ܕ�hT�ɱ_{�V��h���׋tQ�@[�8��Y���.����e,S�G��!�t����A���#�
��>.$������<��$�x��OZ~&�B���(v�uH�V�\�ĽwM[�dW2����©�[ؐu�U�'��4��	`�E=޸���!�D ���} ������^Ի�>����Q��y+�A��2��9���s�%Mĸ�/:�p It)��P�I�!+ F[��gRsz��	�����N���Ʊ�w�ySs[�Y�(%Qex���uQ��H��� �j�6��xH��SA�t��E.K#*�z��F�+8�$`x�}����7\@�y�����H�����k�)�D�]�x.�"q�k\p�nsÈ�����y.��Y8���0r���}��F�`�����:]�!xc��ҍ�d�$��e��=�v�qQNw~�+U"x�.Ss��3U��4w#̭/�ɤcdx�З�ike!��Jm�9�����w�/�#�y��v뷑>�c]��.L$�v��\�u��m�!�\U�������!�v;g(�5��jx�����Z�[��|5R-�З��"D�{�y��v��N=*��;���W3*"kZ��TH_��c<�	�nR|�/Ǵ��T�Zl׭L����rG��A=�zv�"z���}�9s���6˓h}Ե'@�s<�PN	��}:������h�ӿ�+��p�&!��g�W����Z�q�N(t���f����HAz��nbr�aq�+�$���!���*#�����K��$�_� ��oN�,�S��rj��,���X��n��9Z�J;���CY�0�z�(��pj/���V�[=19n�K��WgӾ^�e�����4`E�E��oY���R����/(w�2��U�;K ��Ia���`@�����؟t[���P�҈ p�*>�3[yjό�8
xv���1Ur5p�._�M�o{o���\X���6��)�U��5D]�͗��M��lz��g5�
�/�e��^�zG7���*�"���L?��&�ܭR�|�`<bc�%��_Z������㧰-Ļ��T�a&��M����ްf�r�i���8�v�[H�4�J!���������@^= ϛ�F�r��u��ʬ�$j	��#�LQ��3�S�o�h�N�Po����q/f���	��D��i
c�X��ih�D�$�n����'ޔ��f���xp��������^�S�SQ^�p�9�e��Wc�?U��u") |�ʟ9���e8�@/��V���Rݫ�BN=�8QC�-M-vP�}T�h y��R���`���Wq�h�\�#�ީ
F!u+є�}�6�)�K�_�^�h�'�&�fWJ0r!��� *��ʈ۔�mq���S��k��:��w�LP�v��V�?rN �Z�}V��p��U|
5V���H}ʛh�iu,�F�^u3{�C�S(F/u�_;����J���W6���ψ��xq2�T���J�A�2V���YΌXr.����q�`#�^&|c���{���i"�l�������4(�L뤼k�]|=��rI�%�J�뤸e�}��}��Jљ.g}G�A�с|�{�LC�ﺵ
�"%�O�/n�J�sGk��2�؂Jl�m3�N�6���)�t��*��Q>�hU��.�g��ϥ�(�����������J�0��M|G�����	_[=��yB�_�ujl���iF������+�1lyH±�^br�ۃ�fA�	���lG�խS���RlQٔ~��j�'�������}�q8�3��%���=ߌ�-])���W��4ȗ ]Z`��B$~VD��-�_!��2I��`L��I�[r(zߎS��|��ڋ��\/(��:�eiA�6JJ6�u�mv�_��k�@Lu>��S��-����a����G	�c�n��&�o���X�d��c����4��10��6�s�y�2�]}3�փq�t�C�s��L9 ����7��^ Զ�Q�4�M��#�\�'�0�/�i�*=�OF�EK>t�r�
�5�>6�B�s�l� �Lhg�C�������O[�qݱ�Ҝ�����:��B�r�^���Dz�d4~����q��%�&��zzF�P(�Ia*�1R�B�L���	�p�d="왗7Yh���ˣ�Pj
T"�A������0��5F-�}0�(����Թhp-�T:����U>77W*����FWֲQ<M���&�0��7��b$+Y����||C!f���e��#\G&�l�en���w��|���{+�;�hHi=��XkWf�Kb3���O��D�R�qv��z��Y6,�:4� [��ZW�o}�C��}E@���&㒃�TL���Q4�ӼǙ�ǅE����4�����e�KW�|�#���)������=�l'�� 4���U>Ҍ����i�,X��=�P�P���]�����~vt���[MJ����A��tD�这W`���F�_|���^�X���鿮%��\>	qʾ���w��:
rZ{r'��b0JV��|�}�Ȟ�)Wvc��z��A)+2��iV����1ȚV��`<7R~�KC,8����$��!��#Y�D�%���\\����i���4���~\KC�4Q���$��Li�\̪�
y%8B\:��׌��^���5�������&܇*�Ux�Њ]�?<ٕB�ɪ٘�?��pb��V��d��~���5��S	E�@+`mu��,:�˰W�O�(�  8Sl��2w_�]�X`z�] ��E��6�������oJ�'�B|��@}��%j�V���;Jο��jM�Y�!��_��q�) �f������+2��JOr�2��T5��m�kǁš�,I�I�*)���܀U����G�Ʌ���o��O���\Pr��/"�LaY����Fm2a�#�;��S�>��w��7�a�B砅qd��z�`�,��W
�}^�o�fkb`�>ԽMbd؂���}׃��)�)H��W���21> ���]Q{��?d�@��o��F*P�!��Ƨ�(�"6�|ơ�F���ߵ�F!([E����
�9���N�b��g����`,ݬ�B�6�G�>*�!�Hr�,+nLq?壖�k��
���9~e��P���pbOug���q���oB\�J��>)�-4��@z���"g1������*N�pA��7�$��2Q�,��w^0ڱ8�C��QH����}�w>���Y���B��)��c7���l��UR�}ơ�>��S�j��=M�;�hW|�r�U�t���2c`�r(�)QꟍYn!}�������m�.��|~�f��)�ST�f���F3��������=��I}F\������>>��#71����3�[�F����N�[�G�,KDpdă��)�7)��YL༠���_��-�siґ�58n��r�������hצ�a
���I+n�+�Z�*H�c|����+�)����A4ٍE���x����n�K���v���R���{��%2�:�~ r\���0�ঝ	�<YZ�J���V�~�Ln��r64m�)+�E]CNs�T�-����M+FgKg+��F�5��Z�w�;C�.������<0��<>�'�"�&�"g��F��!��p="
��ն�PJQ�D�_bʥ ����=������r�s�����֨�5O�7@��M������R`�;;���Y4CK�1�H�>@�0�[/��ú�-�ܾ��m�3���rH�e��	5j��K��	8�+ Ԣ�ҟn@G�we��ս'��2����D��k�Л��`&S�%��o�C��!+;}�s�+^bI��)��$dP��Jn��:݀T��BlL�\(����T��ɪ�;@Q�楁��� 9{��Oͽy���d�D���{$�����2��$�)m%x>��E��a�m#�S�|�m~i�,'k�<�_�e� �G����X��d�^�S���
hK�����z-����(�@r������rȢ���"2@1�h��~�h6�����2Ǟm��b(�d�>��6��at�A���%��#Fz��|��Ĉ��q1S�����9c꿂�@�im�z��Zzo�>Q�"�},�Z�L��v���{8���n��3�9�|J48������~�:�U��Gٵ>�O��N�܏�o���u���A+��J*ߡD����p�1(���:c;�N�[���.g!�Dr���H��!L,W-F'��0gx�;>�6���r�M��%Oj]��ߌ��bWm���A�겝 �5��C
��SD�ܸ��K���U�Ȼ�ʖ$M�UZ�&�R����N����G���8d����� ��p���H�Z�),������_X4���ʓ�R��k�a�b�ac�6��������_�����~�t\aJ�1챴?<�&��CkL�?��]J�o2�
%���v�
�q����V���c#��K��Y��LY}���oR\��6�Q�e�=�����t�ut�r����t�4�≢�A�zbK�S�N����L=���T����q5릶�v�uZ��A�8m�e.�j�n����_K��"���Fc�*1�{;($�<V
�HO�Y%]�i�-�<)kmB�* G���'ǉ������O�z�r:�y��!ظ���Y.��;���*՛�U=��j������N�
�%�*�q�L������PP��^d�!�p]��s�_1�L�~Q9;$P&uW�Ô�L�M��/���7�������mW�&3H��$f�!��:�*	��f�12L����ޭ؆��n��1�Q+z.-�����!J�i+]�Fn0$'Xh�S{�:T�,�;x�cq{m��L��M5J�(ؒM�C�sC�-a܊�&��|���:V�-��f��m�k*]��\�Vf�|����L�� �Ɲns\Z�DW}��JyZF�ګp�5�9�s��&�q�
�o�Q��ջ����^p���"��pjBWtT��'���Y�]_�1nx0>��E{I��J�� x�Wo_a�Ts���nN�O1��W<~2�@`�n�T�gO���,cK��bֱ=#�fU�r�it2��܄�@��Zy�:"yCS­�Q�m��S+���ƣ4#w�1(�`h�(�����_f�������m��ޤ�#@�������a����p���a��%��]���r79�y��9���e���U�Q���������v�.�+�O�ͦ66:䵩��[�ْ�Dfx��[?U(���yH7���/KW6���갡w���w�ƪ."U���7��D�d�mn�D��WM��]qc�/���f�bM�U�#��0�-lzL+�V�+3�
��6�����Ơ憛H�	U��_�
�,R=��I�<r2^�������J�z�����5��k�qG)���~�QE��)��'���"���@.�%�0}�N�9����8*��S󏔠��#J�9W���>4�6�[�����qŗ&�����;cS�J���<ѓ�^���R�>�k��TC�d$c}�G����;�v(>zd�Ɠ���m����A��~�u,Bá>�������3m��'��w�� �������6�̞�7B�Q�[gl�;43|�����D��v�a��ӊ��*!�N�W	�[���
�ޙ1(YV&����Ç��伮�
Κ:�M:Z�%f���}Jw;K)3�ʘl�'d�\� ҳ9����k�ĘS��Ē�����N���4a�� $8�9�>m.�<+��z�M�^H�K/\����U�������-��!��ZG��i�'����8;���ts0�`���$Q��x��?�β��ř�?s{(�	�$0=����$�%���ċ��W0+�k��YP�]k+����d�T������t!��c��6���f�SgtK"瀔����V���Wϧ}I8�-�]��҈�'҇۸-��f.�p3�����K��`(+VqO���I��	�\WK�u�S^��_�Ua�~D��[i�	e�U�}j%���s���� <�:7��C���+2ܹ���ؕ:�Lm}��yq)��vkr8�5�D�W�;�s�If��w75�� ���X$嘾�ݼ��/�cu�
LY�7��sҞWt���iX˙�׎�&Z�~���D(��ϨG`�]�U�)f�1��{��;�N{��ڰ�x1���n��$O�����Ekw-��S��B�*dsv�g����+m�b"PU�y� }n�[QB��.9��"�h�r���BM�8��%B���
J�>�oUܞ����<�J�2k�Y�J�i�|5[��e���$��nf�Ғ7^�������d��z�s&�m�kJ�fĲ�둇ae�>M����~�6E�$�q��j����8���n��5�1:pHa�>��$��ج�*��. h�!Lz�s 8?��J�Qq�<�)=�M��bx�!0��C�q�O���I��#�hiJ+�׽�!1����}��@�z��it���.L5,��"�u�XР�R
�� � ����S4]E������TR��fN���r	�ݪ�A��c�0���ǈ =X�!�ްj̽W�!0�d���^9��2x)ݘ���D�J��M�;#1��>�
36��{y,h����15A�_P��!|��D�)9|�m"��6�k�m۾�)dPle�*���-n)g�S�9HgZ��Ť�yL,�6 ��r��{^�IOӉ{6�n�Z�ǩ�$o�%7�\�	����C��S%ݰ����弯e<끥ߪ��"A���Z��B?��u�3K����[Q�x��]�S�=������������#9`Kg���w��#����Y|+��籷����a�=�%��p�#�dګ���5%xu%nv_�J�:�ކ;���н"B�t�r�%��>e1��9hm��8���7�g1fUy��\�l�#8���{����b�{-��G-���Š�B	�<�璳�+y�f����q?�M�Shl���`z��#�.��*}� ���gl�y3 (e�#��b�b:�	H�<r^ڣ;�	�Y�kMkά�
�E����9��y-����K��W�~��ȇ������T����p��i�e��T����(�����;�Ń�v��g�N����n�y5����O�-���cM���Z@����S�)\Q�����R�κG����#@cۢ��eۈt{�#0���Oo� [�?߾�}��w�����x�&1���ɺY�6k���P�,�tΗħ�QmK����p��T�v4�}�y�{c�s�Mx[W~����.�0J�� ��>�5�:�$ ގH����z�DC�c�o���ST�C<�]�=d�����lN؎C�v@�s�Eer�po�Dl3AH�
3*TH <y� �6S�Eb�}l�(P�''x�m_ U��U���8��,;H�;E^�I���S=�=DZ�g�n�Ds��^	F��
/ܻ�����n�(Q���s��Q�U �/�#�n��Lܿ9Lv��6��`(^�W6-�J+t�~�	F�.[�����.̞�K��I���,�*E�����u�I��Ш̕�����<>��B�}��!�b
��^)|�y�55�����Sk\���kʯ�uWZӧR��+�S������=Ma<�?J�������t�k�jf��-��x^���p#+-�p�fkH/��+�Z�z���٧����q�]Au�}]�w־�}b�����ĂcW�e�Յ',�����=Ut� �;��+�c �ٱ�jeaͨ���e�"����@/����'L��Q���픨?��uA�U����I+�����}4����j��BL�oq�ߥ��,����P,���B��=�[�����(���H�v3�����J�#b;�����N<�Q���p��t��%��n��W�L��	���R�8���lrNk|>�������F5]�}`CI�0�j�LL�ic�K[JnrҦ�uPUj�a��Oke8�'rN�#lX�?\����B�-�:yS�g� ��?�N��d�����u�ϗ��0ގm��x2����I���Y�Q�kk�2�\6��ڂ���~���^ߠ�	U�-Z�3�1�m��@���@����b'�l���=�+�mS����2�aY��PЛ�DokM�V�'��?s~�`Lom2���Y��AH[f�4�;�b�*O�bh��]�5w�"�ǕY�Fl�h� �ž(c~j�d�aH!��J4�S"���$���k<7e:�l�p���ƻPRת+��?>�v�.��C�z��.�**�KF��>?%��� �b$�5}��gܖT�TVD�| $�4�H�1"@2[/��	�Y������?�C� V�V:�i���A���t�zM �Bs/�xi�8{�4��p?��Rv�L:٭�v���ދ�kT1d}t��o�m�I����Kқ\���8~�Ch��:�3gFw�<8Ѱ�_�{���b�>��)��)9�
�	�M+fq�@����|dE��M1��[I�ǐ�־��}(�7Y��]�{�fk���ܯKv�3J�q"��#��%b6b���W��MQ�T9�Tz��Q��z�ø<s-x�Eʤ۵�9��|b�t�����ĒF��Ł�͟�w� �u?]Nue�J`]d��_������v�}����2��!�9	/��'��M����iee�Ȯ�5U9��H;ݧ��N��Q#M����T�"?\���ͯ�q�zt�º)�=�gL_m�)�%���u�����=��`�j��6&��DT��`{��G��⪻����=d��@��i���n���A�2��6��c}#YcmG��"���	��kJ�M���# 4l���?� $$5|� jsF�:��0�j.�l�?�4'�**�����Y��f���$���-��W�m�}�0T̼��
�L=A��V�\�$8�c�����r���@T�Jqbeqǈ�es~�@�Q�׭�3��	n��M1s�țp���h�[�lL���=�A"[�^I2*Dy
��/gJ u�h���� �fT�6��2�P��nyG���Դr8n"Wv�*x�O	�x��� e3���?g�>���e	��:3Z�����8I� 7����6�Yު��d)��K[�/PoT������F<˸�^�}�:�~h�g�3&�$uՐ�L)�D�����?�C��1�2���4=�xɪ�v����qwuF�/}p�?9���KS��Y�oт���g`���6�q��S �Ff�T��̭=;��o��n�d�s�X�][�9íن���ZhV���n����]1q��v��U$V>���%�aF�������h2F!(�0��1�|�C��Z&�M�����W�0ah�s�0��#������0�;�0�gMCm�*璫p2SmN�%E�	����F˛�},��˙�Q�93uL3�c�j�ۆ3/-�@��%�:�"��㛘�g�r3��J�����p8��[�96h'�|�??^��B
�z��Q���RˀFO�k)�AE�d�D�Mcsa���n �􊎪�Z�y��HP��s#Cֿ������G0�����.��r��c>�mI��Vz�|�r�R�hf$�����/%֍���N8B���ZK�c� t./@9��
X�/��SF��'y����#+۾Zv2X93s�0Dy��������V��Y�Ʋx��R�&{y�	1��Y��������<�_Ao�cKb��迡�:�44�a=��	��9ԕ������c��^��:�*^6�Ί&k������eǍ�m ���?F�U�d>wv��+��'���q�?k��N¡���s"�cr�mW�\J��Z����ҟA4�9L�*�]$}b���k���#�����p'P>j�w���K+4Z�1��6曂��`���$�<�	4���c���J��K3ޏ���'e�[�*tw�0��x���#���`*�"�iU�w4Uv�k�D���$^����7���c���jw�!�]���������;}P�T)���l��M|�� N��#CR,y�Vg��W ~��w��is��� �_��bak��	%��'�D�B�
0<�F.)HGw��!%��o�Yc���eE�z�d��u�o���_�3�3��u ��X�Z�sG�����,������j2N�E!�8/;��A�^Cfy�0�;4��\!s��:W�Jd;�b�����y%�����ʍ��o����;X-�I�MP+�bQ��'��nڼ�X���`ӷ�����h �Z�{$�#��Y�]�����)��ѹ��Ʒv6�z�A����Tc*�؅����$ޕ>2mw�F���3�6ӜZ'�e�1=1�/�r�o�#��*Dq��:8��U�?��l��C?7W�'r�M�a�b���!O׷�Z�9*���yI���#��16���xcb�c6e�m:�-bd^�a�B�(0����m2"z7���d��=.����V�an�h�28��<��
�kd,B	�s�@��mf�υJ.��gR��+��U� ��,QZ�	��r�{��Y��885gI�Ӛw�NvR}���2]��4׈\ �T��i�<�4����� �e搒dǁ�ï�ٜ���'V�8�ߧt8�P�ˠ�s���G�C�������n}m8��Ǉ�3 ����E�B9�&|@��(�B��)�84.�W;J���!�t���,@#ma<�g�6H*20jn�I����KI�g�=!#,%6>���,��>���eV�
��U�<��N�
��2��ZF\e#�DY܆s��TuHΆ�^���H�K�t�`'�@��r���>(q+_�Ѽ
2�`��9�t���/�-�@�IY$;�_I�
,�w^���]o������T�-��\6�2G��>A����8�*�x�i%����C��,QH���s"-�����SC���Қ�&��F��,o����g%�"�fFsP�3�J.^��C�XFC~ǘp�>ha�۲e6�8�mN��1MS�[�9G|�f��P[���j�>�k�,��H�����"��L$���y5��������:�8F���=�']��XQИ��=-9y���!L���@t��m�Ԭ2���S�!;a>S`Z�����.;\�2�����y�
�|��;�ѹe���Q#6l��q�_A����m�])?�@���@?6��t�D|���@�i[m9��lU�4�I=�8*��	�:�v= s7��Z��9n��;�7�'���Bs3zk�%U�β~�7#��E��ߴ�@^���<�^�Y���V�7�ϗ��¾�D���	,_�fW�d����&d�0~�t�Xe��i^�W�)��Oq �����8,
�7�A٨0��+?H�CL�L�V�?�)w�eD�,�Q{�F��
�0�Gi
���v��pc�!�ɠ�R���.VI2�)^8��e���J�M�!
���6
�? j���q��$��z�υV$7��c&:��R�s�%ȷy�]�#�[�O,�X@��,6�mpB@���$;�O�#2�P�rhr���*��O������jcd�$a�~���~9b��)^�(�M��J�.2l/�&�����D`J
��\�%�������
���Y>����}	�C&%b
�Ϧn�䄢�z�cd�c���q%��7�!����\�+�[��uZ�%7t�@����C&��"*X�Qs�Iάo �A���#mI{3�X��kT�*d�kV;�6�G[��E���n��O�x[(�XG�he�az��!����z8�ej
2#;H�Rd��
kM>�R�T&��2�1u-�GO@����V�73(�T3+���U%V9� ��,K�5$d'L��a�P�z�"�]"�v���;
�	Ws�JL�]ꍀ��Y�f�*\�-�|���{���P�48|ApL����1xk�8��M��6��!���<�}a*3��D�\c�~�碌o��DSsrwL}U(���C0۵��H�j��T�)������D/�nV�?��s��2�]Rk������ �}��x�=�����|bɟ�R?�a��U���$�
|˾o�R����3���!$��q|<nK�嘹*L��\�}ل�T�N���V������:�M��I8B���Zr��b����8&H�4W�SA����\���HbQGG�rk�:�7��c)?���������@b:�<d�WQ��J8�:K���Qic��{�Q���=msEnQ���z��wO�>c�ܸfn��
b����f>�ܶ���c.�vk� ��_;v~��w+qE�'�OA��&���JN��$����M�à����e&�eV��F8���nV`s�@�sw���������63eL)'G� b�� [�6}5-���W���o�[ ����M*���ػ���Y��~��]�h�;���~��YVI��٘H�k�g�0�%�-n��L�pz���ֱ��}#}�% ̈dz���������N��RA�,T���9�A���]�XlZ�k~P6X�'��[� 7"P�RZS�5��tw����c�i/$@���<���>lX#U;����Sl�J�1��i�h��Lu/�@� 3$�-�jȔ��b x�ٹ?����/��Ѽ f�����a�sE�������;N��R��a/Y�
�t/IPmp�@�����,�Sj+~��m�U4��Bz�N�e���3¾ջb�q;���,��gZ �C��H���r<�
��+:��#�@.pβ+�rܺ�B����/Q���08;��tװ���]3_���kϛ�<Be��t��p8�r�fב��32c�hT[�)#aU���*l���5Z��Q��x�eB�	Іg�U�
Tr�/UT���K��f1���T�"��"��"F.�޲��!�l�7�H�W3jl)� �E��PF��>'t�Ԡ�Q =[��Y�����N�駠�?ȕ=?7#U�NQ�˽ȝu��p�4�6����r&�;xr��a�𞨤]�j��+���6�U��P.��n�O��CЌ<�O�$q�c���O�ϔҖ󜃀�Ac��4��݃Y�����C��ߦĹ���|�&*�݋��c_�ulڒǦ'��6�t�ɸi�2�ig���ĳa�!���U�q����P��v�^����U�YY�S>��!'39L�]�O�3	<��ݿ�)�j�3���P��=?�郶!VL�ч��.,z¥���l`]V�3��Sޝpޝ7��Z����R׀�Py�7�v�#��{����L�V������vo*:�)��'d��/��[	���q�+u�mN����*�h~�dM"�O[��h��]�x��d��]mkt��$�F$Do7vQfYϿ�(bT�K�@�g֥>��R�������_��sk���^� ��F��Sb�4^���n^��uY�C[��[-�|�#K��;��Z��Z��j�߀�8��X�(�Z��E��n��02��W�%L[�)4��:��H1c�>r��^��S�Ŋ��/H���[
����a�*5_��8ej [�%�Srv��T�����[�ʓ?�O�A�v��Ѿ䕻
q*����3��1�p����D�����a<e3²�gB����/���܄�󎋬�q���i����j�d[���4��J�`�1^� {�@3���4�1��kɫЋ��m���7?��.�a$"� n!��\��K�a��Q�\(���S����^�����H�I2b=1�EL��s��0�ÉY�K"s����Vo-GF�z%s�m �o���#��̽8Q��l �krO}X�P舛��#�n�����O�^��v�΁C�����n+Q8y�k�cI��67���j3�r`�;+�.�KwS�oJ�-j��wG"�k��٥~HJ�y=�&��"&P-�ϬW�4$���f�b��`�'���[�NE'lg��ܗ7V��+��o���$�l�" e�T�luv���AT����[�7�	b֯�v�Oa��q�Y��bXC3莱
bL��.M�Ώ`�潣���n��Ŋa��"�ʘ% 2��|�pt;5���K]}�>.���PIg���QFf����N4�WG��	��F���0�T8y�Qݷ�����%4h=�q�.�{?�B�'q=�BR�7e�G��֚�Iߐ'��
�p�W�� �|�&�x9ɒ����B�Ҥ$*�	s�,�r�����,T�-�0�}��O_+�G.F�Z��yV���U�W��R�#ն7Mjjv�#2F�0���D��^���� H��������`�+�m�gO0]G�Z��إD��� ������y5�n��l�sL�\���Ew{<��!��8�ml��ɉ]�6z�]��N�NG�E^v&
�/��螬Q��.�UŇ�[²V��������'�%8�T$�'��rs�B����}tǏ( L`��p�M��1^	{�����i�����7�,��>(�1��?ج�7�ƳS ��"K�X�G���*��� �[�F���г��O��(F��*0�<�Q�S���ǠR��w�1	�(�>{��c��Z|��	#�-K>M�h+iݫ<4-3��6�,^6?�d�$�Wz��T����H���\M����'��I��}��߂�W�nwV�p\+�	�Ǫe{�jL��='�KW�)���3>f^�6t�
��Dc�ȯ�����V,S�i�bς$���Ef��U �� ��~���*	{�xJZ!�\s��s���"e���F}�)
(��ä���s*qG�~6ކ��b�`�䓏�^�Tu�+c(�^h�c烈p����? ŉ�R�����U �� ['V��o)��%�%�&�}��b�@@q;?�}��=��B��#'�c���| SeFw���/��R�6vSv��Uj�{R�T�¼�i�˅�TF��˂�������}|����P��n�Bٯ/(�
�$��'�ysv��p���5�Xf�{���D��0&##B%J���4H��d�*�Q���tI� �})c��&��oM���mrp*׎�Ȩ�Y����
>��xk�ӽ��px�x�R�ɒ�g�v����K-V�t��>�rB�rG���k̾ɝ���L9���N���#^6���<�h��el�hJ�b>�.C��	Ԑަc�|H�9�9�G�Ƚ�'	��U��)#��K��xlG;�/"֐���W\0�ǫ�������x��J�'����`gPB^����5y��pEa��	���ۿ�ϰ�z��Qy^�,7��B짍�&���])�m&y+=�F�jR�Z�?L8.�b-�n>�!^?_��	����������Y��M�Zb�}'�o�\�%�M
�(�:A���ףN��<A�+wvu������H�I&ЋrJpl)-�N�鵃�C�-�[�q����#��Uh:pQq��س]� BW�*=������6�w������V�=&ڦS$�NQ��z��c�ߕ�pҫg���|����������$5Yҩ�E�l��K��`_5��, .tpNހETW��780���Aڝ�@{���R�
c�I,د"]񆚗v^+�
:\���*Q��?6���T"Ϳ�X��/m�g,(��g Q��Q{�ᚐW�W]j����AQ�h�AP��7�B�*F(��D�$��.er'�&��J�2�Q=�dߺfZ�J������JW�#���A7�1�H��"��ZV5�:E��M]ze�"��n��ɗ�v�L�1��:VM�"�>�|��҉�R�:����4ӱ�o5��W�z��#��hI�@͏�:&i�OY
[x�-y�{n�dg�{��+�P��ȵ���5y�5��S4Xb	X��j�@����<�'�Lb��L��i��l㐉��ůEM���1��Bp�-�zMjY�� �!M�RH*@��'��z��"��a���d�D�8��J�:ҥ��F��ݯh�3�E��d�U�R�l��BE�f�m�S+�r��?&|3�ե������Uk>	`���!֪��� 2�Z�~+2��rV�hUWI�^�3����a�%>�w����M*yًm��(�{�������ػ<�~���Cjf�&�V̭�#P�@F�����sz�>��W��ظ�U
�����[����Ӏ
���l$�IS�_��-\���D��*�YF ��{/i��+ʫ�S���!@ӺMp�~{�	��$�G��)���<����}���e��>k.Ji�-7�3e7嶨>�P?��-~5`�o]��0D3���E�B�@+��ً�Όgu? �:;���<�(�i�b���i��<���ʌG���GF7b)�h��Ab�ܹw�,��Ԁ(@�Ԫ�p���iYY"�rj{{�t#�n�d"�%tN�Ik�	��jO�`�=�%�c�s�������K]���.1{����57R��j�+����$m�;�Dԗ=gR �0�[G/X!9��¨��{��I����锫<No7�0ݳw� �4���C�a����y�J�Y<-�d�EZ)}�+D(uE��$	��+�w�rb��B�gG9�', ���%q	�Na_x��>����s-��M�u��j���'��1K��*d�0�㞪�"F#�`K�(1���8�?T�mr��v-.E�Q�UVGʚ�L���j����]=�L���K@�9(�u.E㚻�������	f�u'/���Rk��8*pn�!V/5����O��� �F��l��a��������ӹ=�v���7�����F7"d��>~�ʌG�"���Ɣ����.$��.��bƎ��Y�fȒ)*�SCzP�b�-�&�B�8���)��i���ϊ6R�zb�5b�m��Vܮ��,�o��D��H����:��7��n���q9�3P����3U>�W�z$r�iq6�Ѿ(P<t}��
�K)7�SX���[L��qB9eY����R-��)F[�9������l�k��a��JFd������l�^_��{r�	o�2T�Ǣ�d<$��_sT�1W¼L/�����. f5���+Q�ӳ�v踺����n����:9}#������zt�Q���*�eq�&Ռ����A�#��9?��3�}X�h+/�����W��
}n陆.Wavh+p�_�
Z1A�H�ŋE·-ۋ橃�SX��|����ٷ�\�rW��g|�*c?1�� x*��[soUQu�Tm�O�2%���	cxn�c� h��๐��U�O���R,�t����ć[����Z��	��=e��e�2���� iXİ�֙+�1�v�&J�]�P{��"n=�|��ۨ�� c,}��j�ƌ]>���ʦ�7�H�\w��U�`ؓ8��ܛ�U�۩lj���xl��vRh����	
��q@�3t_�l�����U�D�ؖ��Z��EÆ�qf2�
�c!���ך�o,P�bɷnk�J��c�5hS�t7����?-o���P/��ƞ��by�C���IW*'w��^�s�,�>�V��QDU�p�%*{H�>�gg"S�*���;w(ǝ��	6�Ia����3Fo��1lò�bKU��tY��5,}3 z��w��bW=\��U�o�1M?�4B�I�:a�D�34q4n����V���-$7-�>ݳ ��}( �UrΒhz�m/z��1r�kX�� �X����� �=��nOnhfy�날��c�>�%.j�3���j�s�ˮ�&o"i��u�zb��BJ��Z{�����T)^#�� �ZOF\�\C���xЋHwT��v@�= ��z�u�R�#t13aG},�$��[$��ǿ��-��Ъ��e�t��X���V�0_J�3M DW�~W�5����jBї��'�K^�a����-�dgm�`} �L�6�=�5���(�(a�B�c���ki[箒,�8��-#~%�#�����������'��*��a�Y��e�
R�l|'���RQj$�H$$�����4\牖}eM��C�Z�#LX��Mro��7P���R�M/��� ��_�����QY��v�!zH��\��NN��F3BM^�(�|�K&#.w*��5���c�Ͽ�mLR���)��o�'��ft :6�����k���J���!�FYeyc�^]�,)�ܛ�˥�-�ԓ����N"~b����Ĺۧƣ[��Tw�úhD�	>�2J�O@��&��?_���.#�#ne&'�=�� =��@C���~@�C��mޤ�4�d����)�C<<u���{s���o����.��Vy_�yg�pm)*wO��t�ի��cw|�%"��Eq5�P�
�v�9s���v�[�35Ә������0Z_<)�*���_T�|�ϗ	{B5H� .iW,���f������M��ߚ�baqk}�H�[
���g��b�+�j�.ڌ��Y�X�/�bE@�w�5z���>�m�ө#�����²3pC�)��%�a矣��z^�b�"X�b��"����:�Zn��}հ�EHK�S�͈��q�!s&By�=��O�p���
<bk��ɳ8����Z�
y�a2��i��c7�~�Saa-L�6m�Y��E։Q� b3�S��J��g2�x��)͕�r3V�� V�<�DJ��3y}����)LL��6����?[t��|L�����p �K��bJ[E��lK2B�̆�, p����G�?Yr�@��*'4Km������b۹nH��^���w�yc��[���-<�h�����?ut�����`BX!>��m�2�����;�h��;�5�P�Mh ������4����nT���ґ�oVvS�r�ٚ�{�o��OLLψ����� Z�ʚ6V�#�Uq_�$ȍ�x)M���K�x��L_���>z�P��l�B�PܥI5�< ���ٛ� V�2KDJ��lK�����0eS�bn�mԅpaM��W��s�$ ڱG�X6��~6+��*bv�� /&,�4E���:�j9�^�����p�
k�u_�N`��?�5ǬAU��%�S�
h��p��=������~�!����f���S�M��Û� f!_e<Ksd=�J���8b����pzf���;��.OA���	kw$)����3��s׷]�G�2�x�2�5�9.� J��	?�3�Wc�]0���g�F?)Sh�NRD��de\���G Х)x��pYW�1���V�S?�T֌K�������Wcih���������D�c����q�ƹ���,�
�gW#�(�EMJ��;�YH1(_O4�\-�΃����n!�U�EĨ650�r3@h��d��`p�4�Ί[2�k���Oِ�x5�y�_�{#������ɢ������Z����i�T��8ƞ�{Y�1v�T��Ő7F� k�J�D����x�^�\cN/l� ܍��uJι��+R�\�(��V�^W!=C��(]�����"�m�)�T$;r٫�N��H7�8m�P�+$L��Jp�Ny�
'�m� �jη	��W����l�wR�z!��jޤ�d�.��v�&:E���A�`Z�l�=�����9
�x��
���K͐��Cw��て;�R���S�AGO�-H\�X�F�,�Kc���%���ꫣ��e��;�inF�+q]��Ox��ly\��U�
�7?�&F�cS�����* E�f�zT��
����z����1���$a{}�ϐ��c�./#z{�]X�GŽ��<	*Y!��i�^�$筦��u�Q�m�I,?��zکf2�]��$��A��Da}��S"t4m������e@�hKٖ#�(|"<5�ME�v�� �t�������M��RWf;T1@�!�G��c:�*�êB{[��h�Ͽ�y��o 9��n)��3��b���^qE��1�SI�{]E
�������%8�
c�a��4-�w�]m7�fEm��M=4׎%|*f���u;�^��07M�J:���y;ޥ\ܲ��q�� �W���W���v��� ���e ���n�މ�&�	Ң#��u��}w����TT�/m��Wc?�a@z��7��,Fr��1ĵ��7�!T�sJIx�U�&�6��^S���Jm� \�����Č�Gmc[~�����0��4H���A�����2�O��{�e���2��D����ܿ�2����o���������R�CZ`f�2�)�uQ��}E^��
J��e��!WV���ڙ�,���"�s�������լ b[�6��S`�e)�����BW� a������n{2NN�"�8&�!��Ѻ�6˼z�,]�~�:�1��\O��eL�d6q0�I�(�F>L�UZv�*�֡�I5��s��ʾը�n�.0���ACF�^����&_�&�w&�����qȖ��S��c���\�jskL�h(�O�՞��Kރ�ތ�	���7AB����rͥ�*��t���+(�A�.�5q.&��r�Ej*u_9ݧ��N9}�*P�݀�AJg��q+}�D���_#���H'�B�*,'�<_�#���(����;�^��a�kZ�ĉ��:J��#C�@�,\T��;�t��Xn�u�2:�J	�Lo$��`Zi�.��ʽ�r�p���+ì��Fe�z>%�þ!?#�;��q(�&ƥ����p;�'��ƣC� c��y��2}ٿK	�����#��$XN��%��P˒]fV��~�Z�a��EN?)^�>��㵠�u�ifx���A�
t�3�{֜���RIT�ˆ�V�I/O0��Q��8�g �CO�?�9�)Z������靝<��T� Qs�mz������SnE�����{.=3p�מ��7C��?�0bd��-�,l_E[���St#tC?�6�moP�	�::Ӿ|o�k4��_Z���ȍ@�xo��Q�#m+�'ux�3�[�������"��uԬ�8v�+�kԔ�E��Q��%sE��@��:��k�[�0�m��?���z��h^u����ۭ�Y�4dT�! I1���BX���[���}8�%V��y��0�4��%L�r"`��\*J}Yq�`\Dc~��:�ඦ�-���W��G�]�'Rp�>��	�}��EJ5Ikm��l�v�{��������o9<W��Ħ|\E��Q̠�֢������b�#��SP��V��3���� �x�-/��X.�o�>/{I���CzF�+/wbѕQ=��[�H^�׀�Bca4J�H�P�y]��B��� &7�c���է�y|��H��+X;�5��Wq�֬���B@Yj�Yw�;�,�pY<� L��}A�3��8/�׬mA��"g��'P�K�)J$�H� ���L�
|үU�N����<0fqՓ,$-yɠc���o�XUɫ�� v`�Z(�5����l�=�D�֛Pĥ�,h�`ox��%J�&�E*�H��P�	�\
3�Et���b�$�����`A��g�U;p�D"�`��d�0�y��}�.Pd�#�Hj/�Xa|ꬒ�\�dW���A�ڷ���@	#:]餏>@���}��W8%�
��#DљFv�|攡^�?��@8�~��&�\��[zH�P����G9�DW\�"����H�#�&��g؇���q��_ݦcBJ�4���^�#��}��Ë���k�Cx�6��'gE���7���&��a�l���]!|I�إ����o���E� ��Jl���y.���;>X�G�jt�s��g�����g*q4x��"J8�G���/�]��$��V6�����|�:�ه�_#E�s]�Ru��ui5Vs�&=߬0{�f��Q�h`��G|�u01�;������F��qtƩc�X���NQ�8�<�Baɑ+@}��5��O���gj��s�'��Se_�Z��)D/b7�(Qk�<�	�$��$�ڔ��PIp��������a�u,�|8�� �KE�3��^Jsh"AQ��.�:�t틾��صӤ������0�R�C��9m���.̌�zb�ӫ���/bG�Wp>[������TZ'-�
���qɍ~n��!Ÿ��*J��I�zŨ�׋�#�����G&������cT�=L2�y�,5�w8zOed�ἅkrp*Zh����l;�?��Z�ة��N3��\�Gi�xG�zR�y��b�5�=�]Ќd����9W��s�ցཕ��+��N�O��~�=���8���۔�xx/'�s�`؜Uu�:�u�y�Vn������hwp�[�#&����5�Cbғ���p��y�ퟴ����A��l�;��?��j��P3�X-�Ib��Q\I����&���O�9�4��MһRJ9jG���8�a��Jdi��Pu�]������WcHK�d�{8�Mn���x�"#����x��.3�R��L��#/k�(b�E
�������m�਱p#�'�iu�{6�v�"������]��wC�R�B�grId�|�R5��x�}j����*9��d�P�����G�j��n�@Ct�u`��/��$-��Ϥ�����ƚx�
���F�}��ο��NWe�!��SK�o<	���U��k���M��0"�%��@<�5Oj8H^k�����َR�������P��Nk1~}���ޜ�G�k+�֭_��Dm�����e�z�Ъ�0�	'�b\of�~EWް���id��H��ºCgj���#�fC�I�^V.+�+*4屻�p)W� p��h�xC�.Z��R�=-��2,��c�M�0� ik��T��}n$l���d��)=�
�,T��ٻ��PÓ��~�k#8��[�zio�4�����|H��jk��@�I��3�ǵ��݌��D����p�oi�j^�1Z��n�Ǡ=����'@O�S�>����6�i���^�z�B�uX��Ɲ +*F�p����(dᥴ��*}���g�����M[��n�����^�ƹ#+в@�e/_�%+EJ/|��|�_F5ş� ��k.�n�"".z�
�I�JuKj-	�[�N��v��)��;ҚRWƿR��RR9�,��H��:+S�G���,�����1��uř�<3k��bMm��a߰�='*��3� �M�w�c�ɚz�I=6�=TJ��q>��'wb�m��\#����C�j	S�N��w�)���;+,2h1�v�EZ���_�V�<w��;�B�yF��$�ۡ�{%%��n|����n12�
@x�
�a0�T�&�/aw���뵧��%��!0xk��b�>�ջ�b�\/-��)	_q�%�D�X��rΘ��#�������/:��n�d���$�C��6И�b�N��hX�+uZ�M��f��
�����;�'-;���'�0 ��=�E��>S��!�ݏT���;��VF׮���m�`TV� �U �
~!j�R?%�{���]/}�c���[V����O
k�3ڂ�1��_	�͉�n��jyA��[��!q���A�vS�N��ݍ��J�,���:0N|�恇Öl��[�{g��?�Tn�=/f��DʆZsU���z����v���I,,m�z���de�q# *+ʎ~m�FJ�{]p������O��=.�}D%ݫ5����8��_���YN6]��M���k�S��P�+��~��`��C@�XL�~��#ߟ;�5��\��G�J�Yv��	�u��M+�ߴ& ��!��X�ފP<z����P�����s�{�_J~�L��r+]tT)�4+-l<�~\�*>�.��/�`g\KH+N��!�S�ѡ5$熰���;�G��+��~8ϻ_���c7�{#L>����Y@�	U?P��G#Ov��߻��KYz���rPm��,�v_��+��@���4�m��^�T(l����,��sizvC{獇w,qI�uul�4Ӡc�R�ҫ\2���ޫdxC�);BX*-�����#�j�"��a�C�t�m���ʱS����Nݻ�h��I��WX��/j�ͣ:�[�$�O��d�UEu�z��\��2���\��Q�>���.��E<�#�"��7��W�� ��#S�ðY�p%��:��4��Ҿkt��M�D�"·�z�Q 7C�Z���ƚ?�쪆18)!>Mc6��
��-��	DC���c��_��q�=���`���i7⿂x%!�\�I 3���N5~���;Ώ�
�X�$��7l�;� }:�����������������y+;�ĩp�a
�%����M�T�w,�h&f���5�����$1 ��/��A"fr����|���j.�N��<���~d&�\��d^�X���b�����쪜w:�d�K�1���k�J�0x�e(}�e�.]@d�p!�J�u
dR��Q ��ֱW���t#(�dl�_����ba�Fd@����/���k���K�*�+����l�)���|�N}MQ[4O��$���0�u@��sO)�Kɽ ���oa=v����9�&�.(6�+�6J�N:n�=�DyGHܫ�rU9�ε_yQ��7�$�ނ���>��O��9����!��"�5�Sɟ���s��c�zb�"�״����x�Zt7�0E��
��0��e@"�L���b��G���i-Qc���=!�-��@ݾ�Y}�;+
�ơ�%쥿J��:O3�n���Kˇ�mW<�܃��� �yXQY^,���>�������f�7�"^�^+��2&�E���F��F����q�0�w�e(�0,|}�����L��+g�[����|�*�eL�$�{� vF̩��8ԋ�������Ymm������q�i��%>���E��y.�߁A?m�2����4iQ�_�28�ɟ�-�,d�S�#�;T�����қ��X�L�M�7Ȅ.�������Xk&��/� �ʧ�_�7�5w��B��/`ŌgE�������%�z/�}���C^$v#�ʒ�W��Ѩ�l��?'Ҋ�g@�v�~�Y\fW,��W���Հ�Z���'.=���J*�Yy/:m�S{
;tQ���g���V����T,Y.K$;^/F�7e6/�i@=�l
��#�n�����98�c���D�7*HA�Ơ�V��xd�-�z��֭�]��|�_�2:	%T��?4��b$�_����J������v5�KC�2�\�W��C���V�5|i)iB����+V�Yf=�A-n�|ʫ����Si{[6��m~9��e��H<��V;O�	ٳ�OǬ��(-Vο�	z�~f�MP�AL�O�OeF���4;��	�@UС��fY�V�N�<R�6ȗ#Uu*_G�E��
hi-�/"�ŶKs{
�~�5�t�'���G������K�O��&������!ޕs��Eb�Vÿ�,$d���j�h�.��U���o+��jߗdj����g��E"��
;({OAG}�FC2�2mqN&� ���y�*��`�c9I���\6����1��	S>���Y��-L������#g���uB��9>�����^1̎:ާ��s���)���n!:�7Ȼ�X�R�:��P�6�֔�S��|��&야(6%��9R)¹ؽPw��]
L�������4�Pj�DY�!H�r !.,�F���}|���X��� �F�����U�+���k<>.��'�В>���؇����Ƃ���<��5�*�<�'k��DbW\�b���r�KQ)n(���Y��>��ƴ��� pS��˪��|���XAy�aE�lk�V�����$��Ϲ�<�D�N�[X�K��D�	�Ν��fK���s7ZP�K�*uU�'J��2�S�ާ�pNC�h<�,� y�1C{��A���|σh=fu��v�
�h�K�Q�W�8�[\��aHD��_�x/�9Y���0���̨�l��̔�oho�Zׇ^ˠ1;�ޠ7����[EӺ&�Z�v���%��f5,�E���:|>7
w� r�����Ub�Ӄ�#zb�e��n���P��-E��Q�JDڇS��U�\Xಟ�qy���7刷ZY��O��ETX���9�E�:zp�p?�v}�E��7����3��'�i�Xͳ��扳��z�c�ƐQx�4�5��V�kd��ĸ�o\|�r�B��f;�i^�H?P���YRߨ����i^4f̫�Ő�	ΛQy��MӌI�� �d��5.ҕ40����%I]t�7�}j� "���(�&�->���_Y��q�f�A�P�$ڨ'�����@|�����pp��p���$:�C@��M,�v�|�U�h+H���*�����0)�� Q��8V��,�C��`���YPp�)԰����n���#�Nɼֻ�"���e�2���X����[Y�QBN$e�1�b�d\���
�8��\5x��o�Ì��@_��`5�����!Ys�Z�1�w� W8��	�s���='.�j��p�]*��/7��DN߀Ҹ\�Ç�:���؋�^_?��2�^ۆ��ʦ�W����a�gl�DPv�S��'o�]���L�P�����ޑV����V\9�0��9��;q��}|���L���ĳ-� X4*������L�*0,�(HH����F�����۱��qp���:Q������H���A�Zn-��į�7N�\�/�F�:���	�y8�[l.ͳ�����+U�����������	��"�S�t�~�d9R�+wq��^vZ�pQe�����TT��u���0�J~�O	�'�Z���_�)/�{z���|6G��w�2T���c�i"+��3�@d��&��?5�·BwB�.�ZӤ�=u�"�'ǔ����������"�
J��ň]�o�*�č'H^���Z�<#$�E}�6K�%���H��Qmo���\�n7V]x�Q�i���`�.~��p����>k�_L�)[��7p�{EK���-ӄLu43N�o6�.�F �uړ����2�{��Vof��WG`$'�E�#Q5�~E���	���ځ�>�]�Op�����P�����5�J�d[�;�f�c�ò�0���LX��ߤ
���V�������`Ũ�Wm�7'�t���V��*��6i�G%f�(�˓���F��A,�a��>���+�y��F�w��Z�)��m)j�� ���;��)�6���xG]�N+��U�̓vi,�5����e��Θ!?�-t:G\�sy@-��=�.��� =r����k��s5~ZOP�s��X!��q���k�sk����-� ��(c�bйa�J(��'�F�~�t�O@I�}d]Y��]m�AŞ�-$Z�z2������P����E'�]�O�qh�gdvReMW������Q���I&n�ËP��P�7*� �:��;�9»&���*H�	^���t[�kR�T�?�ׂ�-�#J�:F�F�{��5:�����~�d�)
�
����� Η�Q_�����pZ�Z�n���b"�duA��I�(��V���%�rH�C"@��NK=���v=�갓8��Xx[k6k%��B�r����%�q?��`��&5�g?���6%}e_E��nK]��WYG�Z���I{�R98 }�yn���vfl���mG�nK�}�Q**l�d �N }y���O�:���A>��0�(�J[T^�e�K�^�=xo��Z�?(�+�����2�5�4��&\`��Ϲ/K;|�N֜��е�aC�к{Nf4l~[���
d���Y�"�;��D�̞�L��M��l���~|��d��<����U����@m�xWP���SC�aGǘ�V�h�W����0��\�Fs��@�O�}N��ƭ�3���$�?���s����a�^�C�ǟ�P��{z`}1�TG-������qT2S�cf<��c����i�G��h�w<�{p����XdW���G�q�6p��$t��~f鯃��gU�u_������f$0
TX� �;����@�L�H��he`�pG������ʨ/�-K��܊7�q�M$u�f���v�,k�Q�u¡����nvȏ�*�^������e�i�L�U�d�Mhl^�pU���x��qѦm~��`T�������R-�X���Hӽ��]c�m?[C��ْm2�t�՚���DH��_�^c��.�Cq���zF
s
�4J�`4�$�7��lņ��6��&4����DQ^����R���=���5��"֖�u���m���6
w��eBi�b��׍Z����Q�e��Oo-�:V�>�.`_jׇ�*F�T0���ON�~���A�3<�&�d�ԓYj�:��/0���G`>$׉)�H�����Vc���9�p�O9B�
wISh�Q��ЇԔ��*�K�a��4�����d�[�͡�ǻ�&6nY�uV�+ѐ�(�Q���H��Z�Fǥt��
��_�2�M��g�e�ח��]�hB�rV�%��[�w1%;z�]������H�d�#��بd�L��[v( �k�i� �<���1XC���|A[̒�}C���:���`<��,�->-o�N?�D�hr5x�{��F�O�W�̘���n-��_�bo5��3��?��'H1u-�S̀���;a��yb���L�Bi"�����}�iP�<�B�fNK�]�����b�RiQ~3�?_9aZ]l����
=�L~=DP@��1U��\i��%��.w�u$9�.���ٺ��/�C�0�=��Y�e<�/���l--��U��~
;��ח�a�Ȁ��)�ʚ���"��(�l��kp��������B���zG���F�9Y�v(�J�Ƿ�JTY���^�s�4͒Đ�t�E�Ί�	XC|_���X���yn�Z�tM@�Z�i� �W&y#�w猏��J:���Jh��-�� �p�@�\S�D/�F%�Y�#�
��3w��i�\wK�
�|��k�f��w�%aߓ(7���np{k�ʧw�lj	��k��՘vx`8!�yv=��V���|��G߫.d1���^ufA�hEB7a_ O
�8�e#c������-<�:A�
�����Hz�r!{��{�J��-�#��X �OD��D��,��><��q|��s�O#��j�$dT�$�{FV���ї�z���l�Д,�8)�-����c�����d�6~��$	�y\W�57:���m����!Z+J ��sJ
�4��a�(�re�Ou�� �U	��8R!p
q����`�nsC�
�A�G �T�)T`�9�|*�|>�?2��>�g���~8Έ��d%�fڷ@��Q����/��� y4[
@c"��G�-/�K�2�3םvUT3fX����PP�X��[h�b��T��ͩ�������3�> ��1=J��_���t�7K�<���I%�-�q���� ������#��q-�7�%�lZ�}��I����.ǡ�C�+���3�=�8x���2ƻ���U��V]i�'?ၐS�p�2p�N]�v�d��P[䳬\�M�o�����+�
&
tq��E��L��e2��DX��Ns��%����4Wn��!o�Io�z2����E0�Z�+���3COBM��z��V��?:UV�*�l�0�'�/�`�o�Z/�������~4Va�;X<|7�r�ܢ���d`19]dh�0P�2B�س��惣���E�F܁m�͌���~d&�>����1�B�a�u��穗�z�4-@g���Xx��r��g��S¦H����l�B�#R�F%ć<��o��֟n
����l�𭥻�����mS$�!i�~6�B�[p���ǜnu�O���[����[�n�:�8D�*d̓f�O��,�"��]�zD̮�t�,$F�?�90y��H>e���.��{�����V`Y�ă�O��X0��:���[�&�Y_'��ik�)鄮s�
�w`ͪ쓥�y��?o�s��.�7�%"���M�B��Z������q�Z���9��&�{����4��MS�6�2�j��;��
3ည⦞�iX;*�������&-�/9��n�@.G�s���1�������Wp����"�3#�Ӷ��M��	$�����k�� �x%�������,����H�Hm8%�U��i)6��K�D���B�殍㉩�7���K���B�>�a��H���&����e�1�h��N�{_��\�H���y�^B0�H������a��"Gj��ww���7�Z�/�d�>�!�Vz���,���f�[ê�=�[m:��
U��̵6q� 4�d����K�-D��>7�3=�X�ϥb�/����J�Z���n��Q0�9P��.rN�7k��֞j�u�.��TOI��S[�4�D
�~R����"�Ѐ��rҞN�2_8�`�uyŸ��X��l�`�#(!��Ҫ���f�+��XS��*Q��*�G��+nS��B��Cli)��9܂Mi=���cۊ�Ǵ��ItQ#Ъ>��A��2��FX�9%�]�<���>C���z�&��6�Ek�	U��!ؽ.j��L�4�;%����(a�2	�B����3�&Cɩie����,]�(���O[�(��tR�W(������ν55��ڎ/T��z*�q��岍�����U���Jz*Z�u��x+����/�Q&�A���T$����<�JS�l΅�2�m2Hj%�=��ʟ~�J��n;y4��4ݬ����d�{�\�%�ى�U���>��eb� ����Ԓj�����#)�G�T�=NE���Ahͩ�<r��6�BZ� �^\�~����Z��h��e�:����å<�-ұ�[[F�\���b��q�=Po5#7��91��Q<�Ib���8�9O~k�\]��0�l�1�^_��xY*f�@�#z̠ʯ?x��+g��3QZ��b�|���f�%+B�IA)���#�L&dI����Q������k����2�k�1j��%����$�E�J��6QT�C7+�>P�,Z�WQ�v����D׍ר7�Z}ΗhFǁ��hk��
��dD[V����^�� �h�"�Vkk���az�6�\�4A���H�D?Ʊ߭2�x�%i���˵b�`����YÆ3�(�޳�SW�,����5�MhzCe��ʔ23R��
PH-#i&�u} ��U�Ho4�V8 V��G�nS�����1��F'�b�	�^�U�0�h�,��;��ؖ2A����s��45����EN�2*ϰP��r>�������b{������b�Ud�N���H�oz}҂ѬD?�h7�0�w��b�ؠ�6AeO��h�+�I�����o���F�0߽�ٜQ�ǋ�2�(��k�aIa~Q��_LG������ʨ�]�����-Q*P?Q~*�GDs-���������}2ߜ>$\;�<;od8��ѱ&��0Г3V�&7D�9E�
�Z'�0�fZQ_��H��� ���U"YP.����<����/�9M���tC��L�fN�vkl%�6�2\��9`)�4'>X<b�<J�Ud�>�49`�Q-ޤ�Šznݶ���a���~ھ�19�ѣ�z��W� �8��x�P��	��DK���]HBx��Ki`��xn��=����$�?�!z�RaG�1zR�ԞM��$R_'�S��&+�^9¹�ĬP[�VJ�:�Z?�ax/�r`�O�f�L�����A�'w&��bb}�"����3�S�]W/Q-D굺� ��\E�MFy<��nA�w{��>Z>T��ZrQ�6�0�p�`� �;�|�O9��D� �-�����	sRG�Ȣ>���dC�(�A�9Tq���D�C-����m�Nc}~��[���5D��3c�Q��_m�������g^*���>�*%����*����>�^ =+¥xUm�$�-Y%��8��v��1�ƴ�&X��a�*�����{�<���Ot	�0�� ��t䕁�e�~B��e��@2�d����`���
(�Bw�P�G�͖��~N���_��{
V�Kٳ%��:|��k-ɓ�ͱ�6���0� �n|H�s���By�pp���1W0f�P�f{��ȯ��9�6I�G���Q��TvJk4�w�u0�@&�s����� �+�ǲ�3�Z3.�$����t-F�4�cG�1�(�g^z�$�s2:V�[��K�	:V�AG���Ƙm�(k�)��dL�H���L|m�,:g����s��"~�v�#]Qz���®c�{\�d�����6�� �%��͟\��SZ��(�A��d9YRv����)L�O"����oɟN|#y��ǆGƛn����d,żR� �{��@�ʲ=��,�ExQ���I��3^�ѭMy_Q�P�i1�Ω�B���ٗ���(�-�&��3X!��C�5���WkWY�<���㍚����8d��۲�6��>�=0Z���W�>���#�g��	{FW��7��Ʉ\+��Y��0v��t��zm݋�	�:[/�Uk��^Y��WŊr��lAt�
�1T�TfS���1pN�%`E�d;�=��j�ƭ��:ME���V��"_X�:��95_��T�� y-}�}<���	ݤ��Div���d�-�"�R�$:�9�6��%F\��O�,�#�{���|�3r�<�1s|Eb6
~O/ϘL%��U$ʥxe3E�9w������S�^_�y����;�,�=II�I+a�0p)�.UG�G���r���ל!F:	���혦�F�}8��ꦁq�]-.��doZI�]��%��Hݹ"�M{���xD�9yV}N��Ֆ�����BL�MP�aw���=a��e�����#h�5;W��<\R��i���>���̯#k�A��W���"wm~Jq�!.����T(����T��~&%�y�����:H��X�	���a�Q�yO�	�
M��0�7��g[����n��G�Z�.�@4��o5]T��j���bkE;�����;�f�����9/}��n �ȜĔP3Q֖����سl�O�@��T{���\Tn$��!n�:nZ[�y)D��t�B��bTQ55�1���c���.�k�槈�X�Rn�b��*��=������K`u(`�xv�K�65:O��R�}h~|�����
��l�y���u�`0���K�{�� JKYLs����/���x�����P}ٻ���Xn/`�6Rùr�LHK{h�j������t��n[���>����]�������ŏG,��(�Ӡ{��|t8p�7A�@\�n2�m�ږ昫�b��>��ɐ�P"�g"zo�<2s��k�t��D���krT5���:	pR%�[�87�U�2�ٗ	X��<ZFY��9� ��ߣ���R\��2b�}'.���O����ɏ)d���:@�N0�˨������tQ��j@���Ğ�1$�HͿ<��:��E���y��7�}b����,��%��0���4q��m�*��(��z������3iD�K��h�g�e@�C=���[�a��
0���ϕAD�2�&(���tп���/m��6ea'����ާ?пu�Ằ�{{[&��{����2��3�p�3�D�?�)2|���t)w��-VRiϜ��-Xҭ�����Kc8$][p�� ��x��cCo�.릻�W��Z,��2�L�`1�؉I:5J0r�;�u:OW���_���G�dKq>��񣀲�UTQI�ɤ�4B���"�s���}T�hȁ '	=�q�c4|��a�k�d�M�/rF�sV�[��4�T,}[z_&�od$$��9��j����:��h@W������pe�u�e�p��9�c�Se��~-*��L-Mߙ��{�r���6��pw�a9�;�&b�ZA��GDΜ��K򶞛���R'�����J��Ƽ ���ڤ�`�_����Q��/j�G`b�M�v�g�Tc���h1���E�`7w��vb�Jl��W%i~~]^:����Y�ԕ_JM�E�l�!��?r;�ҢyU�i�W�mإd�5�e�A�%�~�uZ�e�	�o��Z�GJ8ё��� �>W�^Ae
\G�M�04He5���$�Uwsg,��z ����cx���Ǝ?29]j+b�,�ʙ���?�X����XiΡ{�lm�k�B��iTJ�f��ǫ�<�<�2��qE}���;�R���
8��|�)A"	B�q��mJ� nܐ�%!�S!~!��(�b%�R�@'X�@��H�c�mA5&�ʓk���R�z��܏ib���4���|��X}F����,�?��K���rVgb(���%�`�,���ߥ�.0��4�������_Ռ�����?t�9���[4u{��2�0R�i{L����B��[��	ǃL���Xd�6<݀�GX��WR��*���#��� �51�ws/�Z���_�_���W:x��J�����X�m���X�3�]�\�~���Z����".�иe�l�m���\�'~)q�G�'*�fb��!��i/�/��Uʚ�҃/�Fa�ߖ�[���̻���+�1�����B��v�H�
��O��t�v_7]�lO�"HH�u ���|u'��4j�z�6�_��n �^4�]��?W���Ҵ0׽�������,UKNc7�%4��|ir�9�r'm_����Γ�-�<��'�!�o,g�3W�`.��pښ8��TJ��^��pTk+�Kq{WHOO�>PUC�����*��N�;�ُ�e� ��w�yeUqᆡ��͂-_N{2Z�;̧�̍����,���ZY���E��z�n�[.�|��G������>�[�&���Nj_�Ø�D*�9B��ޘ��/+�]#����N%�L#��7�$��l�G����R,���g�l�E��0D�w���O����{�Iՠ�UJ��ˠu� �Y ���Έ�b�����O���N d�1�P]ی9�w��䛡l �n���S�R^��c����_j �a�ϩ^��cL���	]i�W�s	A��v��</:m�)�4�����2�j%���lJ&�~����ܒ�����q�ۑ0���0;��G�z�ZQr־���<� �3�5<�0�B�_��$D��*�=�آ{7���=tڧ��\ �Kl�/��ʌ�%eѲ�p������$�g��	mN��'7P�ʃ��W���@� �6H�!��,�Z53�6�������#�H_�l��_��mTh��f]Q\���I<�N�-���L#?�T�)ʨ�!��Z'�l�ʅ��ޕ� �_`M(ݎ�\�Al��ͥIeϾb�4WM#G���Rw�Ϝ+��b��|�<l�ɚ-�̀(��O���,�b���5��:4��2$cY��l��@��6H�3��}Lu�y,�@6T�jgچ-�[1<�P�z�������(�%-�-"k�<�Q���ܩ�0�z�bݠ�T�]��5M���岍��)k���qh%u��	f�	\\`��x���.�4I���CJME�3�.��ǅ� ��7�P�3�޲e��)Ln��F%��k� L�fr���d��5���aNN���Z~G������&n���f���pҕ�љ.746���8@1�Xx�o���h��y��x�`�DP�ь��Dn�lǶ	�}������<H����2��?�].�<sꏢE��2��8�%�k��4�%�r�?1�ک����1'w*0Dޛ:�{���/�Kose�����8:���-��T�!Ρ����-�%����{��'ZU\(E �L�=��]d�G�^��2s�8,XmI12L�r��op�_o*�fD)a`�8�����b�ʕV<H8{�%iYew387M�2 ~�w�C-WL�Z���Fk��<f����5/<@V�x=S����Z�T��h�Z���˽N�LĊ�Ae�����/7A�et`�)�%�l&b�O\�U�����@�Ͳ�g��E+Տ'L,Wi��Э�|�`���"��O�Y�IP����aR1� �"ǟ��l�1�-v��*]��@��y���n#{ٓ
�c������w����[w�b����Щ�#Ń����^`�K^ͤ@��μP��"��L�!���(v�;�}��1��d˻��A���a-�/F`���#����5����ћ�.@U��P��i9$~�n��|"ky{����1����H�~f�z��v��p�� �C�H��󑠃Y������-ȋ��'x�K����9X�lC���84&��Zy���.���}���m,�u
~ŰP��2����T0V����n7���Fq�>�Rd���2w��d)A�H�ć����8U*U��r
vpК��O��|asc�J ����tr��>@�:�O�?V�A�����8@Y�I�Q|�B�?ۓ�\�"�+P�R5r~
�U�n�Fq�3a|�1 �|18���>W�(cM�5fUpx�{.h!Ơ�B�>T)Sy�	��l����+'v���T����͎��=3A���qK�6��멙cH�D��t�6k?
�@���j�ȇ Ż6��/#��T��x����ig8a��&�;-WF��� 5$c�+�hj)t�V�M�˴klJ��䁅��3C�ގ��d=����D���:�R(yS����x, Ä�|������~�;�M	�FE`����M��*&��^*�{RC71��V�$��s�U^�;����'�I��M���|)�96��1?����uw�r�H��Mv5T���kLf��V)N~I�?��Չ��a�I�G5�2�م�B�C�HӔ:5���J�����]����C�u��טq�UاŧtIpB�����J��6^咢d�����|ԓ�-� "��>�U��p�~@������\�bbL��@&7<�7��J�
������B�����ݳ4ֽcph�,V���8�����@�������V j2�LD1	'0�`�<:�'07���@�:��)���'�����(��4�5��3�gd�����Z����U�۰�D�h˚�Cӡ~`:�\���=f��>��6ꡜu��/�"��p�g��;.�D����t�O�$���Əʙ�NdǨj���(��8����"���t%�+�s��	�ӴƮ*~����}]�ݘy�β	�x�ƻ1��S��W�V�B��Ƙ��04�mv�Pfj�����r�<�E\���>�Q����#>�O���`�i\R��|�e�=��D V��\��4�����_�*��>l��*ڝ�שc��@fx5����@�Ė����G�G&�;Q��� �yt�O�w�E�Z��߆���	��E@��jEcRg����R��Dn�E_�t�X�����=o�"���F�^u�Mu�h�d:���[�It$b=��4�h)�9����7_>Y:wɣ�.�5P���84v����^�	�hG��Z$�23�Ӝe��G�%��y8�?�����8��~���x�J]_�:�z����E&ЈK	TżT�eI�����Y��~�Yh��f��j��	m���,Uаm�$��R��J���!�9EaɱEY.���`D��꽱/�p����L�l���`[�c`��ܺ{i�:,�e=�O�XC���|���a�*|SAyϓ�������hخ�I�zpGh�06C.�ګ����c �pK�WM�{!@5N��a��2C�~��D�Z��5IzՓ[�fV�v�:%�Y�m��vG]�L�&�W_�	�UWh�I������.��xP���Q:d�~�?gl���p����H��`jRwu�#�����Pk�����fm��GJ,�\.��ޯ���i��d���9k�r��+3c"����u�9\����7D�pR.Xt�i�OP��RX8���\Y3�v��аh�k��˿��Xa���q�C�[���3���'|���wl5��|_(=8��uù��<;BI�Fe�Z���(�b��������ȼ�SVs�xW�s�#N��ߠ&�MU��tIX!z�&�i���߃ܢ�N�%���8��e����P	�v�B��թ����`�/����^F�9����K�1!ܗ @b��,=>$R�`����o$�}��/��IS7��� /5�����V��$ ��_��>�A��a���!z!.M{�6)";�Rc��-���mDl˭�5���zA.}^r�X���Eua5�(�j<Y�#�R��`q�%i� ��
��D��F��w�h������$b��b��m��OL,'*?�����b#�L:s�A�hӽl?/-����	�OC!k���Í���7
�HtMek�M2����P_Z�
z~ 7ld���f'�/X��Y��."��o��Q14c�jޒ"�X�[j6�;�N���"���l�,�6c��~l�.��P,��ƞ���g�r��1h��Ņ���6�e ���[���Q4�xp�f7}�1A `����lE\QL ��r0ɍ(޷���+�MY�B�h�3�j����@v;��J�S����zDj�s�s�9 �4-���)��628�3�D�,X=�
A2�U햁�h����Je����\D��2�H��	�^	�#C��h^x\�>��7����b{ǝ5q������5�N(/�&��Ŋ~��z&x���E���O���Q���䉁��`=���$^��5a&�?�e5���{���ܳ����m��N�t������ 07��E�UJ?�BLJs�ͫ��&�)m;JY%�>��x���C}ˍJ��OO<�I".�]IkDA>��լ�lZ�l5�o� :�:�`h^W���o�����s���w$�ؙ��QQ�
R�H���`�������B5U���	-Z�7�޾��7��l���*;]k������/#E�S4�&+�G�CEP�_�ww��1[�e`a����Y��π2Do�"��֑��ˉ��-M<�]�s܃�.J�w��DL������c>
��Rt�s@4P>�-�+8�?����8�6��R�W��N�A: ��~:0�B��H����@s�3��䎦��P�R7@:���
�w7����U����B�č����|~h~9ir�uZ�Hm_�U�Q)��6bhB�j��N����Eg��^��i�8�ׂ�߸�{��QYl!���+F����/�DCby8L�MXh���������8�
����y�h�i�<um�����m�/$ mS��d|�����*5N�k�-���t���Y�2�-`�_�`�|g\~2�g:�j�kD}@�0����P1��_M�a����Yq1�d�g2��	W�d���n�Q�i�ÞgJ������ʆ���U�/�ֆ��y՟���fM�@�ʨ�ÑbX�)W����
\�Z����d�F�`��������T9���Aە��r�T'k�2W�Ns�]a��-�ۊ��
�������&��iX��0N���jм�"JLn��0���m.)N?5���ŭ�g���"؆J��OPj͊D[����P��L�Ev�2L���Ym�|hA��S�^v��o��ah��~ XV�|�K524��+��#�+�(����"j��1]fK�_��};tI���j@?c?����=aH;(���� �|��rHu�\�SM0�}@��$'��@�u�i/��ͼT�Gi��3����g���u��d�X�D�G�����0�j�*�^<���)��7v�����B�^�%c���8�[�2�R�+����,z��L��I(�£@�s�u
7rE��1o�{�,���˚Q�$][�pCC
�yP�ڴ����LP��t iȩA@��S��YNh =Ì\�����z��u���w�,Tz�@��41�pc�9��a�h�CE�lj_84����Ͽq3$�N�^V�h��<�ULx���IrM�~)f���)��U����!����W掅êJ~|���p�jqF���@� ?��|c�9w�:�)����{ȓ��Ne��"sC�v�����"C�-ؚz��N��7)���C鑝\�����񢟸i�HB� wnu���t��7��J۾�ΗvNj>]a'�P�(���<��9
��'Ƹvv�$�B/:�F.�����P���5h�ŊA���fj�*�g����s	�~�+ow�c�$���\���B��t��;^�a���~�"��s�0���̦k��be��䕬0��� �yNC��i�!�0Q������^��q4�>���s�0���Y�lTB�Fb�uߋ�7�Q�)�w���D��ј���v�X�@7X�C�r�0�(�(V'���`�C}+��k����������eෑ�bg`��g���P,�9�1"j�$�v����霂��!��_��>�3Ivat��Sw
��C�P/I�3έz��`�V��5������j�����*6J0���]	�$��q�߃�����|u;�A ��<Ow�X[�g#A���\�rG��y~g@"����n �-�4Ov~P�Y9������ =�LP�Al+�h��Z�G PU��.~&����up�W��d{�6�S\�2�0eX�Q؃r9fnJd%6ĥ�)	?�*�z�4��`����c\  �V���&��ι�B�v��lj�D�D� �U�i V[Gԭ�ǉBOEq�R��v����/^���"�I�m�q���{�����R ��b$x�L-En�����4��'&6p��Q��[Y��W��^���d���m�Q����~%U���7����p~&�O�T������C�W5�T��G4v��͚��>���e�2BQ_EhK�Ȕ��Wu�O�7)_ţ!���7���z_�k��_��#�}"Z]���2�|v��e�>�L@`J�̎�ZZs�M������ʅ�E 4N�L]떌�y Gr�	��������	�aL�eUN��B|ܿ=��3#@���	 &��p�5[VW��	�Q��5����|+v�T��C1�{�?"�&?9��hZX�;�'��DУK�IG�^*�$ʤ��/��F�0\'��|+�W��L�:C�������$*��o�1��O�c�o9���]���J��q��Ϫ�͂��d�쳩����ʤ��Lc�{��8�	ˏ4�_���.�J�K9��D7O��l�>�j��$�ƌ�Z��yb�n�?�ؖ�k5��+��{pd�D�q����c�/r�G��*};��kP��C�.FҤ �,p�{4Wr�ꢉ���D%|���(T�q����ChY�T�ᆴ��e��X�k�PeCL�^{	
�� L�\2m��,T5uCI�M�1��$��d��~ѳ�bM��%QD蟇-��l`[�K]����pQ�2 �������]�ZU�[��Bעݪ+ю���ۿ�h�"B�ƯҦ�8����8���α�Z���;�h<I$52�/k6�?2��%kLk���	���h\�[�K��l�R�\Ҳ�/�,�ymK����D$�-�}�����Q��|ŉO�����D�7mx�X1�+qi���5��=�zQ(*�n�gg޻��zD&b��*�f}�7Ԝr�$��l��K���m��ӽTb(N2q����^ݳ�:���.P��7&9�.�g!5����y=�wўY��0_�1����s[�}
a^lQ��.�/�QѼV�L���BQ䃏��3�kE�>�at/�,I:R'��:�OQ�c�� {���h�䂲n��ޗ��7T>X�4������p�����q�8Iw��z��?2k�
�1���UM�X+�0g�@����Ka�1�R �S	`��a[�[%�H7�fJ��b�R���v@:N��Ӧ%�b�g�H�b��lT�d'��m��u�u�|�{�{�Ȧ0���Ŵ/��n��Y����
��Bƕ�
g#�$n�@t�r$Ď�Niz�aZd!�R��(���:̗ n�G!�����G0�@&!�{�z�ם`��GF3��Е5b[\�L]�0��Q���r9Z�!ޏ���\��58���=�.����H�C.5u�����<��n���i��1wܸV�B����^�cy�"`�wy�;{-�����|�K�oi߲c�.���U�)�&�ˏs@�=�1~����#���v�s|�{{L[ҟ����Ć���Ȧ�;!�lZ�� �Ϣu�'�<�+5��Y�cԆ�S�<KXȳ��4T[�B"��k ��ԅ�]M�S����2C?Z�<�yYєsq��-�Z��hyH2�9HJzQ�j=r�+�0�h��[��g���gn�C�T3h�3�I�N��}�7=��n���T�_�V�u�|��S%{��c���w�{�Z�zK�w>B�πﺽ�}*g��	�5�oDw]��m#�H�X�ۗ^L*�㞑j�F�X�[�T�3/����Et��	��(Я���7��B�Q ��j��������~��ɮ�6as<i�31��G�D� �ꜥ��ɩ��,.����5�@�o?�A~���{�`�'��y���cp�c���t����D_��s呿�;5�����K�AB�S6I\үz���>,��uh��TN�<XU��8n�mfg(TwA�CV��u�p?��e3��I*��p���:��>�>3.M��%�>p.�hp���d�y1���y
f`Ae�&	n1�nV�QC�4i$��M����w���s��	�oM�BT�P��f�1H=	nŮu@�����xR���Vr�vb�p@���%����z�PCw�3�jT%X{����پC|�%�sdc��>8H��y�yW�� |ČK@�Mhu*�[ÿ�!\kX*�J(�V�׉+����S��}\f|�ńo��/�î������_��҂`+�0��H��EAc���#���)C�5Ŭ���qM��"᧘���E���]���h+��4�F;�[_���{��j��ٵ9�*���k�$���ػػ�c' K$�#�.&�����t<��趚�ǎA1����PI�B��O�m�dO���@so#$Wr�b�ޒ��G�ʘ����-�eϨ�e^��E�qOh�æ\�`������+�23�J�� ��]��j@�_H�������Ht�M�W��Pq�z�+=�
��'+=@|`3�c�Q ט���������n�(a7��̟��E�%
¡�:͆���@yM�W�h�3�XG9��wK�1y9|ț�~���Q�SW��T�}
��D�O���s�����?C��v��Q����X(I�O5������@�5mC��	**���i�볜D(�;ha³Ws*y-"�M����fDKx��9eZG����*X$�|w�x��R����qv��1×ÄݵF�-�,��p��k�jȍ��]�A���Y�ژb4��м��r����h�������8皁��$¥6��E��R�\98�ʻ���?�����|b�&|���2��ēa #�+2y�����G�0�+ۓ-=���(�
�Mv�ucO7���nk�����;Q�5	<�)�c�^M��؀�4e����W>�n��������aI��l/(n��pK�YH��K�?im7xy��vR|-��Ś�ķs��"is(�2r��u�gr����h欆�:��CN�.{P��Z���ű�UB<�4�f��ب���O^ߤIՒ�U��*KeW!�ZH�����˄v5��64_e;8�d~ԺVL�Fُ�J��!	�/FA!��p[���v.r7�,A�CHܸT~Vw�]�Y��F�b/�[!1�x�F�F٢/���m�I��wS����Z�_<�a��6Օ�U8�KU̎����;NoU�z{���d���#ֻH���զ�ٳd؛�U���X�c�Py@Wܡ�ڃ�Θ�Zo��db���Kҵ��ud=�78��%n��4��˾v����~�Nzǭ`�c�[b�������B�^�Ե}�����.�2���KR�J3�@�pmp[���.��j0�`��p ȝ��ܡ�9�B��77ߺ����q�97�#�i+�Bw#q�wӺ�iS3�ړ��bR���O\��ý��V������1`^����5-cP3�E�DN}�Y��/Ww	Z��_B��{��!q���[������SN�h&�*�0/���S4=+$"�l#*D�@j?}S9�7/�m��/��kfpTc���ܺ��A^������HK^څ�3��Aˌ;d�b�K�g�i�:��?T�����]�k��֏��U�M��c^\��)䅊Y���\�����%V_d�ɜ�DD� YEY�*s��ί��>���eci�V�96�Sxh��z�L�g�`�q��`�M�h`����MCC��J����=�Zhh����!�`�����8��#�O^��_��&1�\����n.k3�^fRn���M��.W��F�������[�;L��>��5��&
���M+�N��H�EF,^f�@��"�K����ŗ@��+|�t�!Lj"�R��tNzE�g��}Oa����:X�������cS�`c�T�茻1b0Cٸ`��7)t��ţ���/��66��{���Q�n����=(��-pw�p�����������X-�O�ik�OvQ�B�ek���g��5�p�35<Z̽yy����u�z*��m������s�4r���+���؟���y�ʈ�Q(A�+��J��� �EO>ӯpL� ��/@k��lz^w+�#�U@zSal�m\�U�}�pjF:S�VMh���֥	3���$/Y�^��{I��������2��}&���>8,��:Zp�~V��z\����u���1O;b�J��o��1��_o��Nb����}�ë��g��Vc��rXkL�'�ű��u����S46�cqy�_Ÿ����a^/D&d���:@$��Ͽ�XDq4=BX�ؒ�����T���H�&6�ˡ�A�a)Q���Y҉��ۘ���p>y��e�n���~�����VmT�C���a�U����|���W�����S]6Mo�!F�P���^[�	J�QN���2��H��\?��l��௦!��R[ߪ��K͟�7/�:��W
���L�ɤzU~�����6�
��S���H�W��j�������2�+^�Λ�0�_�~Q)fUz�ֱ�S+N�r҆��Y1��QzM2�
��؍�)�G�gl8�	�焲W�~����\����o�8�a���y��n��sM+(��d8�n�;�:�-��{�x*��G�����6X&��QY<ko���18��yиT�kz�L��0r'���J�Zx0�3�xϗZ�k���X	C�F�=Kcr�] +煮���6Ln@�O�Wn�nS/zBp#&��j��W�B����uEcD��!����N�xe	�b�xEz�ڄ��������W}	��i)H��7�_\^�Hs?��M�	vdt�Ѕ��UE��y�書Խ�g�vH��}s�Yi���2�ڍ��=�nz�酌��X�xSš[^��䟠�����;�ߜ��r��\�Q蝯
~e��om�ښ�>E��;=�d���E{ɥ:���v��ݤ�Rcx~�7*t�Q����j�#l��@�M��:����{��N>�
?,:���QWw�J�HT��Y���	Æ�nz��\7��=��� ���@����
�<�]�<ֻ�OY�E%(���,��Gs!�r+e���Eۂ�v���oo�q/�`����vm_�+V�(!?��p�	l��n}5٦,�Z��z�A@X��ݹ��!����cZ�j[)n�6��=g���L�Q۟�t"4�A6�����);K�9k����C���6���&�܊@�x!Q�D)��?�\��/#�/��)!�V��M��x�]ɴo �Ǿ,[v���������Q)�n���M�?�5��h���>kP�����`^e�@z0��Y�)�,�_�д�h(kb%�VbJ��2w$�(kN��O��ͥ��^2����i�-H}�W8b�%����p7��2?j&��o%� ;>���(�]o+�!�K�Ә�tՅ���<[+{E���ȗH	��hD��s�VJ��.#vH� ½�ξg�߽��k��������O�:��m�^�\�
P���w�@��W�^9�E�<2X1�j#���[�t��~��aRI0�45F��exp����'���0�����0����L�}�u�gi�+�1�WI	�a ��M!�`M�ͧd��V��St�*9\�]���N�
��k��Nu�ۢ�1��)��J�kQŻ?�*��ce�PE����ǟ��9�8�C���?X��xgېI���ܯ������AR������HT9������F�x+���vm��1�?��y 8�8J$���]����K�ЇWf��������N���k�Ω1�\���#�1Ku��@.s���m��a�[�a/pז������p7�NK����*��gQ��&ogɚſ8��qr�2�G�:������A=��o؜��R�>� ������R��+���H�?AK�_ ��������]���������fw	�3%]�bY�0)�>�c��t�
�l��b=p�		E�rI�.��PXϚs$5�:>���c��]���Ӝ:?3�rm����b�vڵ>e��"�d��_�I�K��i����(J�H��>����<o!07�A�<���`xyVP|�3eB�dfa��Tb��8�l2���w�坿�5�J��Y��Du�!�/���_��*e����Y�L�����H�yiS�#�(Z�&5�f�9@�P�i�$^�%1�
�ߕ���o��b�l
�͸E�`���E��N0A}�BX��sS��~,�&'���rX�40�?��_�%���z�v��R%�����T��"�9֞m���B���H��J���5�7�������Cj<+�2�f������š�9���xW	��޼�AC$�p�m����+��F�-R+��O$��Հ��N�?m��PJr}f��{ ���Vf�D�%�ԝ�f�T?�o]jQ�]��	}��l��mU�cW���J9��p�&�("W�t�l�]�7�j0t|�^G&2�9��F-��v� ��|�5mPQ��0^[��K��I��	��ו�0v#WD?�m)��E�60��R55�9��pa?���r��I�ϐ��W[�W�b�?�9�:�F��}-gbi�-��/�w �����J[�p�t��宛n�<z�����K�T����K!!�{����S\��	�<�tI� n��uu} Ɂ����U�_�o�/���=րO�,5`���1��|�ݭf�Uk�1�t�I���� �@�S4��6cmQ7�j�@�b8 >���d+�1G�ԦV���):|�t�.){�������s
��皤���}��|Ed��
�v�-�U��)}�;�����p����a�/0f�֫
^�ۚ��m )Hİ9X�p+�F�$���=�w�PVQ�YfS��`�f����ka�6���+u�F7�p2��qC���|��q�O&t oJ��1슼�8�l�d�[�w�ry<��l�YQv7���؁�cvw͜�L�@B�1>�G��w.6lg}Z(�����I�x����(dHz��sۏ�>�S��ǎ20���MYu��>���������}@>9S��<]����Ѧk��6�g_<�����k�Yȗ�Q��#�.��v�D��aK��0_,Q>X�Y�'Q��Sgs���=v���}{��̑�/��Bt9Oi[�ش��h�?���F|��i�̒��ӑ?�47k�����N01��4��L���0�O���xm& ^�=R1M�};nl��5| �k���X� �<��Ib0Ei�|<o��pyH$���+<hv�a�D � $��d�?z�}��k��O~Yn�P��Dg�K����%a�L���rI�Xk}�[<­��b���eQ$&֢`g�¿�)���2�^���K|���-p`�ol̶ <��{U���QC�D9�Tht����ʅ�)i�$4�$M�e� Fm����SƢ$�Ω�s�����;��|ʹf`����%O}�!f�/f�V���;I��*��r���0䣼P?���V��oi	z����Q?]T�[͕8�'Ì$�ʺ���x��O�!쵽P��T��Iݬ//�5׋�H�'�+�W� ��t�a?u�H'��cr�Ӹ��|���s�$����36�=�.��v0�i��Dլ��k��=Lf���zHqORr��} W�����Tt,+����n����ߚ�V�"���j�dF	0���o�s��cy�x���J%��z2��"c������%8Z.@t:G4WFXuYjw)�qG^<f��\P��+}]���-�! �Ծ��@C�Կ3�B`u��f^�w���lr
?�e��],�p_�Q�e�Q�ۮ0D�_�p�s�Q�]4O���L�n(�0q��h�f��}z��J�3���ܓ�>l��˟�]=�a��Tcr��Ԕ8�U�������Y��jPG�s�P'n��D��IN��bwA`��*$�I�� �:]��,���QK⨢qX-���7��������������7la����ȋ���f��QW�B/�J�WDƢpa�S�����v�_�6,���TZ��D>I��d-��+U��m�a�5�@բ�۶2����f�U+�u����Fo�.�k:tń���$M��bz�2r	,���wV�h+m8;�[�T�M�J�i��>D�Z{���,b��7�T�c��`ކ��I�lD����NNڀ��4f��[Kg�z�Y3=#�Y�+��~��.��®ب���<mv��P'F���Y�X��N�]m����U}�W��`Oh0Vq#�"�9蕠��"x��|���9����� �n�7F����a���8H\��ԥ�{Qk�b�Z�\�e���rsk��F[�j���4����(�m�[�B"�eW��g�x������6�!	��m��x����R�!nT���E����20�y%?��'�� ��R�:� Z��pb�(P*x��$bG�"(��jJ�)�\c�����J(`�z���Y	ག�z��&*xo���f�c�)�}*����3@p��G�'#��[�Ny��+}�\v�|�^1��P�5t��s�%�3�5h�Y_eg'c��1 �E��M?�t?�b�E��Sx�OJ�T���ȭƥ��,���2|pJ�Y8c��6���9�]2�ߦ�n�f����r74�<�s,��̽�:�	
Nj��M$	��&l��a0�Ġ֫�X���{�r	:��Z�{���iSk�f��|��n
kK���j�5��=����bT�4윑2X��S��{�C�٘P�����WC��d�3�<��URF0A�B)�m#�Q���U�o&hj�������j6$�����������N�I�ӊ������w���r%(��att���Z�%%t�⚲d����@V��qf{�v�g�����rK��}�.F�e[�(7�����̯ҡ�UFg,��2<"���Ct�u:i;̦����t(9S%(PM�k�D�����=`_^�-z�L��>���0r����G�ɓ�gB�\�XK�.=��`Z�7���k������Z����,���Κ�+��S#��2>Bϓ�]q�Yٟ���4'�!U�W�-|S�;d���Yc}	l���w<OE�Ai5�t�b':ƙ�StE �xK�sx�������o�oVf���С4����Դ�d^2Y��B��b}]�
}�w�d�]��;ױ[N��ґwB�W�<4������dD2�g��{Av���:���+��7��!���AxrϬ�fdG_�����B�����Ԟ'k+�5�'^�ͻ��`����O����������Q��]�-}��e��7�*���������oH|�i>R ��ɡ�&��ѥ
���N�� ��Al7F�{��g����m����f{qdR%OQ�-[��/T7&�;�l�ŝ)Rg\����G�8�*��D��Li�T�iO�^�g�{ϴ{�"����E���+��b���xJ�v8�F+��U��VOD&�0��j�O��؟�Ƌ?.Z���I�mts2ݜ��v���>�	��/S3�bߓ�Y�@9Ky��鏼�J`FD���#�i��A�f?�
��t� 	҂���v��]���zi�D�YyX���νf9�`�_�4��\�׮��'�	u�h}�Xav�%g���so���-�w�[���	B��&
#(��$�Tp?�Qbe�����t��
G���֬5��������x��	�J����w�bmpI���r��d�)h��T�YX`�,��������:���2�xEĀwEJ�0���ld��$�Y���GWW:�J�T�1w����F�՘R�}�A�<T�i��;�����y��2�jn�]8�I��j�������S�;(�=I<jk7�H&�+K"���H1��V��=BUnx���ښ�m�p�Y}u�@iڬz�X,&e���r�.#������2 Q	��x��0����#��u���y�Z ��̠=Eլ�n��Wʀ�Z).c�	���Uي<�6�9\�,Y��4d���^{ౣ��`BXuI�����uQt�2�I0��cf�y0�}�u�	��6����mb�\9K�7�"�晞P���_�][ht;W5k��|�
@5@��mD��Q�	gu�M���(�Zӊ��x�m��|�˛J�����D�AR_u	�b�$�	F�V�~6で.�R�H!��Y��g�C�K2y6����Փ� U&�돯���Uu�8k�������_�[#.o H���\7aA7IH��1p8֜&:`�Ӷ��0J�͓��f�� YL#BIı�(�lj��Ӧ��F�e���f}+��ӵ��n˘Ƹ��
B��+�Ֆ�����C�[�ӣ+�դ� ?�B5��0ϝ}X� 'CQ��^t��#��/�!|�������R��W5B=���v�֩�|x,�cv��~��m4����Mt�$������R��1��d����J��Qʺց�Z �7V(�L��BV�}���{�$�����Zd�y�
 o���K&�]
C�,���mW���S4K&7�6���0|i�P��@?���u��J\�q&C>n�0E���]�B�9�2�i4�R�Af��]�k�N�6Z#��@�M�{���o���<=��}�)��2{��IMb�M[��$��_L8���`To�F�� m�qz��襏L%��eAZ���Ћܽ��`D�/�L9xH�t
�����R���~��"�ۑ�t`C�_�wī�W$Ł r^8�dp��|euz���1fu�|����ӮK�;#�0������}��)}��ۀkW�`K)J���k��h�ه9Y���W��g�����!�9��ۣZ�z�hr��@bt�P/}]����W1��}әb���x�����C}���j�����k����	���T���qu[4� 0��e1L��L=���u�rA�L������L���f�R{�|��;ı�k����j9Ó������a~��d5��PW����qKw�����z��d��{�v�.FC�1�`�$_�<ҥK1�q�pLS�6�� ٭T��]�7���U�	�;+]w�ȩ��J`e��4p34\ºVC={�����]M���X�@�4�[o>���m����*�rד���D�K�|���ծ;�g�fC,j,hϿ�� ������9	�� �v��imv�	]�#����5�)	k:�\�����(�n�5?:ދ���ʸU؈�����j�D'�(��pO(�J�!���>���k6.`���"(�s +���T�޳�8�A�?��\?T�l��0B��=�A	HaN�
���1 m����p9Ne�cd=v�i��<�ѝ������[�ƺ���^�zI���b%�Y�i���:&�T��vS����sCJk5�M���<��i^ SW����f�X��T�~�	��_��_m�7�=eۊ(��]s�P���*]��F�%��|i�sS��I�p:0��d'�x��Jn��f��P9�GcJ���#�J��U�ӭ5��9o���%�1�N�]��U�E����8�@O�3C�Ç|�Zl�u��v�>�*u�b�;��|���!6$)�8�6a�W1�}�S3�p�P9y�>�H\!uS,��Ѩ�7iW��7�<�F"V���9g�u�*S���x��Ov��;+���!�]�(���F�5#�"��ٶ �\���k�d���P�@p�v�O�}����:�����r�s��0�mt��hx�����U�lȼA���2������X�S�!�#�����]q�Q�Epl�;����-o�^h�#��P��$tb]��׿���3l�A�yn�L�܀��FթD�UM�1�K5���n�L��P���� �]�s̟F���ׄ�#BnA^5Jf!6���;���x�{�@zk�Us}nu�,q�����j��~��|j��%E�
n���0���w�J��|z*���u�4�����w�N��u�W�M����*jWX�����r��������~)�6	�>�F(W�E.Y[�~0F�`���Lx8^�ҵ�)�!,Z����FY�t��L�\#m�2)+ëO�����ޕ�$����^�?��őj�c��c;��A�B<�k�'G�5�+U�_;����׽-ށ��	Kk(T�,�+�_�g�v�[�#ӡ�~�d�H\� yۤ[���w`B�UL��g�F����?̩��R	f��<ʎ�6l�uߍi�'�C�@��I�tY�Ɛ��[�7w��$v�}�Qq��?"^>T9��Q/�M�+��tt�U۠���%���M\�[]/���w���c� m��L��z���*c<"j��c�������t)Z�C*6R���sT~��A�ň#���#py�p��$÷�_��Ւ����&���E���4�	�D�@�E��BKg9�Ĺ���*3k�1�6�>=�z(�����K��Y4̬,��P���?��1�����,�;Pz_�FV�Y��3��Q��-2=7�R$ W1OȆ*�۰S8�����H�C}y���LG�MVa���G�.���ûlڽ*��5q���S����,�r)���C
Ü����Ï(��5y/�[���j��h9a!��8M��P^i��D�ie���������
l�p�WE(���?v.Y�9��4)���'��Տ��&�uCW�����*v��y۩�_�[z$R��%�x���5z�jbe�5������R�|�5�����������o%2����xG�t��X�ԝ�z��"�B�[��6ji1�#�_��&<�.��%��0m��h��� Ҡ�O;�K�-��kΣ�E�!�W~�8qpAU���]���wln���0��w$��i�+Wȯ���]#���>0���[�Τ�%�#�5�v��M��n�J`F�7&��4a���o&2����n�o9�zaY)���6�a x��D7���0=6�w_��(Yax����(����'IuГ�@^4�5	V_}BQ��cSDTx��o���x�u�c����q��P����ǰ��8��J��p�t��Ҝ��6��4��0t����05P�4R�έ��S��L����8�>�� ���ˉ����z[��,�C�����b�2H�{�NK!;=�5�r�Y�G'�,��_����Bax�&��{�o]@+e��"�16V���}Ja,%@��w����e�k��Y�w��R[�5�J�B\g�)Q)�� ��eJ�$F[�`s�:Ol�xb߭l�g.�hk��ߒ\|�X9�WdX��gf��J+g��#���##�A�an�hƖ��.�l���9�\&%���Y�NƑ��d�Y&�=T�����Q��W9|�SK���.��ps �>�kx1��,D�t���=�=�9۸J"־!7��m�ׯ�T����x�C!ss�}q_1 @��s��֭Nߠ>�?.:��,���^��F(��ۑ�Su]��J�@�����}�na]�aG���G��5�C`��)�4�@�1_;{+�B��	n�KB]�&]����PO��z�Y���ikk�:��#1+i�b���( �I�	{N�9�-<QzPl%��hA�(щ������3�d��c�S;��^n��n�|*f�@�ב�XD=�j�w��j[8�2�����Ν��=*��ӱx^^�V��FD�'"���C@�7c����B�1�+����6nrt,��/��u�D�&�s4<����H|Nr�{�'�H�JF�H�o�5c͹SsvZa��1,��t����χ�����{�f�8'��Xe%�r�����{��ܷ�??&xR![?iAM�^��f��2�n�n|�z��m\6?����|dp�R�oY�Y�����0G\�"˟�>]Tj6�_�,�}aj����r� ���g�����0�<fR�WR����Eڳ��?�$_�'�Y.s�����0y����9Q�?��b�' �d�;���ı���zv3�0����V���~����R�X]q/(y�5��ay�L���Ր��=!y�Γ���3��t����
�8���^����~:�<af�'����� �ne-Li4��F�8c%�=ُn: jłv����h
�!Y�j��� �^͝�DM�fB���W�}Rǈ���˄��0�,�:
Մ��	7����6�K@��������Z �r��Y����U�0?D��?�Ā5\�¬o�"B�&���4�oT��9k��L��Qhd�2�L�K�8���U�����xp��rWzH��F�@����m�@�M��_El���n٘	���?Q"Sn���Z۵�{�?�Q�R*|V�Ҽ�c�˱�,�`Q���9u㞨oH�4Ԧ����f�O)Yc�؈x���2�4lz�S������ey�}����	��Mj�!��g�J�*�c"��5�� 6�	G��_ ��{���9�^+���
���Hk��{�i�8N���B)dgG���A�t� �&�",Z�ִ�l}S�K�cK�.dв^���y`�����߰�վ�p�+a�]�'� �����w��0�'E�����h�K��q=���y:�7ID��bi��61�����_�,�/�������>b��V}�Ē��}1Z)H�eb�"P-sv5'��Y��))F��h��Dc�<N�۟�F�rV���<`�J��i#����IA�b�EP���S�AmX�n�J�D�mˍ��0�N{�\c# �vH��b���s
������u* b1�5���\���(�6��o�7z�f�n$v<x�C#͖3q66:|ɦ�ߨ��iP!�fQ§�cFRN�v���C� sdS{dQ�����������}L�7�h ��*�-Q%�4���t��OC�b��"��"�_׾�eퟍ�(��[K
���ݓŜ��,��W��%��	W��	�G���\�;3G�m���v�<glDnE�?�h�ܼ�'�!�kR�X"ˠ�$Z����p��Q��Q�x���|=�~�3
.���
YM��u�Rm���`9�w���0�x?���]�{�Ʋ�!n�PPO3REX���b %gCtFy�ڕ+�GXs�'�C5-� l��L�H�Ao��B��	�arv}�X��Z(]8R�s�z;�?:~g�\.��i�m>F`�'	��8r�[���S��n|���"k��k��L�I�}�>����g��9U9o��}��k��Z���`�v��8J"��H2P��������u�O�ؕ�*� �@K�����2����	ih9�(U1{j�7�yǊ�^��@��6�㮚""�ă�Ԇ�l���uؾ4Z�m$:	(}�r��:d�����z��hgE\Q�@sF��Qp��s�=�	�B__%�`�D )��(x��w��yR����'|MD�I]Q��`+5d���߃zt�JE�J	�3�O�c��@ŮQLL�1�Z�w��h���S��N���샛
Q�\�3"57��Q��a�;w� �z
��v ^�^2�!�GZ]�`��|�����zе5ڜ��j�DW%D����uD�B���컾����c�6X�7<��K��>7�����95����Wc�~��[q9�\d2�nN7�,zR�s��Pw�qc:����p��H��д�Z[�;���8��y:��'���
�(�)[zJ�U:m��.�vy���TA�ߩIO�_eHt��s���E [�2�����Š��X�L��r؊��\A���#FI�	�9�s����ɯ8�� "B�5�%�?��K�S�MԖ`�z�z9fDw�i���(��ۋ䗌��1�7GdhW�qO$v����25U���.�[ w�\|<����I���L1��
?T�����^د��r�������]�	��Hl���j��<u��
i[���gj<�RÇ��A�wɲa��Ol!�mkߡ�.���:~p�O8v3Quj�%����:C*@3"J�lo������UꚒ���.ư����E&�+KMs��i�Wl� �׋[��9�>@ =�κ�����{Օ�w .V#��o�3`����Wñ�Q���Dy�əSXfYiY���*�+Ľ��R�)G�"k�nD�����9�ԫfSW
kӵ�U���>Tw���4�96)���'����K��xd����O�H�ݕ�xT�d����qcU����hg�'o�����ƒv�������x~���P"oq%,�c��hf������<�_��X��k�ߜPGy���-}�N�4��d��l��E���N��!�CK #p%��;�jȲo6�'�\J�e"T�[���ߊxLٝz~^�}��a�C͎#�.?K���E<mG��ȹo��/��=�;xw;�q�U�$��67�¾\��D�Gf|k��@Ms���q�$���*��z)%�A!��z6��l9+�6ʹ���4�����˙b�ýn�oޯ3r��T�s[5|����/WBݯ�3֕ �v%��x�_ԎmX���
͉��������������%�c�:yXg
��o�p�<��t+���G�ZW}���Q1Y�7Q�/��+6	D�p������1\��`fh�E'���N>���*�Ac�"����� ���+���@i@x΁���7����Q�U ;,3�3N#�L��>>"BKZ0�FQ5��W:�b�JFr6��ymYI���++z����2Ѱ�m��w5(�BP;�ײ۠��-o|M����-Bbhz�>���2�vq�(0��J_:��$@y ��W�ґO�W��H�f����@?y�^(�J�t����g_htkp��(����М%�'!�*P�4��q�D�c�"����p�N��F.!ir�M'+�wW&az�A��Wm�oi����7��jn.OюS��Vc�AAװr�?Yt�yF
��I�ēL7�gh�"��>vtpo�%��8ߊ�[\��{V`�v�%�|�Kl�tX]���hL ���0zc�oy�SPK����ĈM���9e{�ą�����yA&�l��Y���v�h��9�6��V{;v�E��@��G~�oQ���H�-c�Y��K����T�E5�`x�[D��`x�,v���?�i4�:�5E�2�F!���tz���U�j���gߏp�k���,��x33/J�
"���"����>C�a_xJ���d��u�_�K��T�S�[Lu*%��Mm��H�{+��z��m�D�����́�:��oo���Z8_�,)�D(�x�j���+�����~2�ζ����lE%��)�nk�H���� _?ő�%3"^8�����o��y��j��)w�@ǒ��;�/�5�,��:�e[�RY��[��?�F�m�~޿��zڄ�Zd��>����?w���7:{Z]��m>���u(G<d�3@�K]����9rffT����}�q3ѳ���ˎĢ��d�4�W�i(���)�S?q�\����
��:�mZ��k&1�$kf�J�^M��P�F#��.�+��� ?�ɍ�\l<�%�DS̋�����7)��&Iէ��.�iR�E̎{�EM�oFƦ
Z��.��}�r���Ԓ�G
F��h&bX��J4��v�c��{�G���v����O�"��,�-�m�ڄ��dcN��F`Y�����Q"���Yd��fi����������@X�\����3Y���_1�l���Z��[�3捚���qE�����ӾD�%/d
��Q��Ye]Σ��
<�m栶�z(m��7�����w��yF��#Y������K�Mr������9�i�m�����zb=����5�>V�������iC�a,Q�F�Im�kE�����z��7��Qy���,nS��z��2��{�)����!��yAx CՖ�O�2&�w����w��~��⯀��v��P��$������#�m'��t�N���x�4A��?�JH ?�O�n�|)G�^�v4؜��O�$�댷�����o/l�`y�V�����g���i��{�����\�ت>̷�4��5�$?"�~��9�]9�sƋ$�L7"�z�;»���h<�`;{��1s-d�E*Q�~���3���@R���n��nC8
��T�`@ e�����0�!�Ol/@�%Ƨ\��U��9wz��͟1M�^������-�jT�鞲��w�M 5�b)>PQ�X=I#2�l�a�[6��\*�b�}:��SQ�L�N��n�� �n���@����V{����R̥�Z���.5�=VJ�D>�Ǿ	��J#�1�k�͔���|AiO�SԦX �YT$9ܙ����Ϫ/"�<# w9��Z� �
D$�e.`?W�K����Z�a2-�x�+�!����ME*|��b����������;5q�|n��*�m�5[�2!���n�v#�%���,|�t�@
�f���xa�w���C!��ĩ��+�Y12|���!���L7��m]�8z��!�j����m��[��%�%m�;0��I�4�J�Ï�ZJ+�i)��e$���*�61�W��˫�Z�^�D�|��C���{�"$^&n�$S��'�U����+(a���z��s�-��>�J��{��#��I�V��Tj�.�?�XZ}4��R��y�1�Liv���X��O��r�*yQ��a!�yx�$�������o1�*��%���oݍ�T^Ce�|��1���;�>��ڃPR$�Ԉ��˗��͋�-��Z�N�P߽=�9�J��>���6b���y�b�o��%\��y��Y=�U�|ւ�1�J� �B��r�.�I�=�6Ƥ��xY������7%�T�F�I+�ц
�b�^h�F�6@�s����R��k�T��#:��$�8؟�z�j�3'�
��sG��P.@����SV����5qRu���g�3�Q�K���y)h�bi�.����G<�5�[H�>l�m�oA�bA@�3#MM4�p��lf𮸡R�ۃ�;��l�9-;W�g��%�G��!t0��rPp��(�I�/=?C�Z\O�a���u����dv��hî�\5h|�W��,oNӮb���Q�/Qj,�X��T4Ҡ���$����ă%���&<�XR�͗:����f���$bQ!y�q[�=��}�:̀䊉��0�x:EO/\T��Zh��qebgy�{�&��8�SM����� M�1����u���=�BSP�ZK%Ƹ��s��7U��w�9ɴ��Mn�����Ca�g�31�}�&��x�x���'"���D��?�
�W���u���O�Ɛ�w�Uߘ���s��r[OD��s_�����U�>��85Zs���l;��q�>��Ie2U� ��4d�
�h7�v$.1���J�m��dz��a9 r2�sk6P��sa���-&Tv�'u�+n��&˫#�q+�>Ic�n�&�qtY�x���:������s/���*��+GH�uJ�ze�UZ��xZ�\*�]R����.��-�{fV[2
ol��s\����$]�+E^�>�f4
��R�C�ŷ�����Нn��g���eº%d�4����̱���{&r!��ou/5Zy=����+�鰅ЫgC9a�w�J_����Mz�8��QF�"5����C�Ng�/Ј)��TؤlT�-3R/b��>OO�;}#ꁷ�v |V)����U��fF�[6YEG�m:C'>S�C(u���B�<�PV%�f�@rz�9��A����]='���G-�!�?�ΐ©|A��"�mu�+��3�����F�<^9��v�m��jl���ř+���H͙�d*��Kn�l�����A�e��5�4��h٬a�{ۣ>XDx�ˮD�N���N�E�u�ҟǏ��T`�5P�P� �#��V^�	���E�VaI�,k`C��>_��d���~u��>�	-yE��z1ߝ*"R:����j�"$�>�az?�=�N���V�����?`L���#hz�32VF*!�?�50��츱5�(��:~#�m����t�JY�8Nn����Q�hT?Fj��	. ܷ}����?H?0�K��(!�ć/��*J��~B!�<��f�����L���κ�|ȣ��L#�D4�2!Zg���#��t|�!>v!�b�k�Ϡ��:�֜ �)3X�#���������K]9ZU�[fd�r_"��&k)��g�Q;���#DnLq��~�{�Uzd�9"�9S���g���K�I��rn��MI3V|��㙎�G60'GqUU2���V��W��N���2�1� ġK�����#O�,������q~�Qus>��|��ކ(�D�ǐ�J�z�_�V�H4��Z9S_Ko���c��r�`ʳب���&�'��$?c�LP�QH~�He
ԩؽ�p�֠�.\�B-��_�.O2���ReȩR��s?�N��%7��H�Ko���l+���[���"j$�wl�(��yn������ז���q��A����:S��B�����~(_:*>��?0턧=,�~O-��
��A�x��r�'V����Z5��C��ۢ�/��?O5msR��q���$Tu��z5:NG��=H���O���x��^ȓ��0M-��;��
(U�t��7�)n{��T��s�&T�y��vY����r��r_�H�
BO>�5�I̫9՜�r/'0[������=�s�^.v���`Ƞ�bO c���MA�Y�pY$�w~ʞ�X�0�G���E�ġhk��?]#N-���fk��>��1�(�hl�#��Q߫V��2Ϳ1���g`��;����Ķ1<K�~�s<��ᐜ�ܞ#d"1��D��}
j��A{��\�#�e�K���Iȱf�&��#�.�9�}6�L��[/�Mc�z�q	2E����[gX9�rW�'g���i `��Β]�*7!Q��#�̱g�h�]�t��I~6=z,"�Q��Vg�5���:��I�\.W��+����*$��8A�����a����)� >�MCu'fU↲����:�k��b|��~��`pXk�����Y ���v��R�D�BDF�e��u��N�����$-�]a6B7_��Y����Xt��4��ꏂ&�EjgJjm{�W�A���� I�4ɚ����Nn��̪ωկs������ڷ�V0ə3ۓ�C���P�A�8U����<�
2�L�/�P;�B,�6t��� ���RP��J�5�,�b_��8d�(�ECM����,I��sz^
k{������`����T+S_@\���(u���!rB-U��q&L�;��̆��D]�ak��<���&�������+��#,�I��Ex���J�:�IqD���^<]@�(��[�d�^o�p���lg J���E��g��?XQ[q��Ay���.�)=�׌b������q�(����I0p�)Oa~}c�T���#�L���.�LfA<{滪�.��k�!1�����G��Cц��%	.��~��x��eV�m��W�˚���-f�����:�C�$ ���/,Sߕ^��<����H{2���DxH K�]���afc2h�b:fv����D�~���g��o��xĸFƋ���WiuNf�h�\��!��ߢ���ɧ��N��i{~@} ����tLZ��_!�Л�P rU�*��8S}��lHo-]D��0��<]���4*����@��UTP>��rF,��Rm��i�|��n$\܋��ܨ�Κ�1�������Uj�MfV7闍k�i�<uS9]1��I)���"-!�d�{���zW1j)O ]kKSJ�WT_fZ�B�k�����iK�o�~� �ص>c��3�V�M({�Rɫ�x)��At{Z�� ��c!'�[b@b6����]��N֟�o�^���d���9�@��{b|o���mS��&����G���fX�AK���iωL�ɳv�I�߶48I�5OEa���"p�/ު���s&T��}�{�q��>�j��=p�0����]���us��k�l���9, �*j��H���~\�	X�	5U#��1*c��$����̸� �@|��{t�C�w�~� %^���Qo���7���灢� ~ڈ�	/L��O��d�x�KPb��D�r��-��V��%�4u '5�s�"ݙ�l!��<�`e`M�{� -O��B9'��`��,7&T3d6V!X�540��#�ɕFט~bp����m�*	���O��(Qy���RW����%)�3e ���?�䖰�z�1fz��2�N06�����#ع�����)��D���)����uN�{%M��::���D���8�R� ��z��6���+���'��W�(+�
'����^[<脵�k��Mm��hu���UO�bp.#H:�����"qNj��&�+�P!�N�q~1��l�-Ի�j'V�Ú��eǕh��P�qb�����y$dn��<ek~!zQ3��J�q�~�^���ʃ�2�˲������I���.`�1�탏��x+�5	�\�א�O��7�!N^n��r3&�.������U%�
���+V�!�M�4Nv"o����y>KHI��?A��H��q��&�j��:R)�:B��\��=1Y-�������6���8TZ�#�H�#�D�,��m=0s97c,�_���S)�Z��f^#��0�d�xƞ���>�8��:V��l�_���I�@�"� ���M�@Y�k�@1YBXnO
��+��1���,��Ln" nB�����s#(F9�]��5���Nwr�$7�FY<w����<��d͵��������->���X��?9�v�hf��B�������-E�$���e���>^_KI�ACj��'���X��na}��9=҉V�!�Kb9��M�g��6�J�䀨=�،��lXfK�l������\ox�_ۘ$�>��ֽɽ�Xޕ�x�(��1C";ww�W�8a~��~��|oG�dP�qk"gd*�����ᒂ�'H�,�O�t��@ԥ9=Cd}�h��b5U�5tS�.���R|���o;�������������C�O�����,���h����������I�34�d����j,���=r+a�i/�VB��m�ph�H���5X�a�\�oA�O�w���46ۜk/u���Ȍ����������8֒�K��N�E~�Ko��*�'{Ҙq,�����.a+.��t���h*r'-u�?���RwPe���i��k5�=�`8�5(�O�)fp��S������5�0ȉHg����ZǛ��!������sd��^ ,P�1�M�є#�EA\�����П�����M��+w�+��##bp!y�e����z�L���h�g[md�2`�"��^�
���⠲��/0�G�����`�;nܶ���N0P�>׸L�w���!���!�be8�K1�W:������(V���l�}-��;m�Q����˷	,5�*�l�����!��O!j�9���U��������u�$e���i�)��PD���g���u������>F3C�i�@+H��4��&�W�`9�k�e���#|�����קH��������n���jK��n��9M�ih�;>��(��<�~���Q:r���]բ/>�4�0I�|�V��
�\mUa����)��]@ �愈0��E��V�Iv�H�yi[�s��l�p�>HD�p1��p?-G��8N<	�y(��H�L�Ѐ�⁪G�7�I5%�d+�����17cO�*ZN��z6��.��&Y/5Ӏr�G	4��jOvlh���I�(|D��Wb�8���2w���.�x4j8�
d&~G���W(ޡ�D�ݴ'�'w���S��1:S��'� �3u�@di��z�5����1˜E]�izV�!�␱��H���ZR��e������h�2o_��A��@ء�mD��9���ef�;k�%[��ς���(bW�W�+��Hi���$��Ā+�#n�e7$������Mf�'��C� F�c�Ya�_^�0(��Z�Ssbd����9 �Paq?�:\]��(�N֗	�^M�L�M��r;�WZ��%�E� �CzW�{���~��%f�)�n�+v�ʭ�y�lIk�U��^c,t$��"��W�r����(p�ͤf!):�������l�ݭj"�`_U�W6���~�u�rb�Y��Sl�Uliϕ{	k�'M[��O@d�TI�7��3:39��u
��V�K�u�	�ٳ?�$��Q����06�S0�h"^I'�;+2OB;��@\y�L*��f��P�bD�r��ig�mi9�w�tRRMea|��{�b�~gהD�O�\��k0����!�ݖ�.��+.y�
����@f��j��ˆk�V����!;�N'��M�`D�lB�=t�RT34��i;�r�wU�`D?�T�o�
�V��
w��!Ѣ��$\�s\��6��ʳqm#�����L:�����F/�З;�$F(���c�Ι: ���?$�M]
�g��U�Q|�N�g)P)l�Q�1�w`;7�o�Ж�M�y��ݏ���c�{�~�11U��K���V��\�+�B�B���&ג6a���,�}�� �ut��l�ܬD��� m%�̈k����K�#�AU�%���V�S��Y�V�}ok�:r�0(3N^����aH�ƀd,I�骍|d��ư� ���k�b�*�i͗I+A��p�*A�%l�aG��1gW����j݉M7y�΅R����1r�Q=G���}����� ����@��ƫ�0--�H�0&#�k�m�
(}�����B�Aפ0ˇ��@¶c�nt��5Qѵ�6ް�C
������n�bl���sT�wT-��Q�@lE���+02ݟwP�d{|�p�|f�.h��~�_9����h�=�3��f�6f��������&�%�Z0��O�ۛva�I�y⣜��i��?C��Z�mc��>a��@~q���Ε<�?��l�	y��[W�"���q�\��XL��*pa���b�!D*nǱ9��q�_�i^4%��}��Z�|��7 M��X�H����B_D�������|'S8���ƻ�GWSyܶ�1��A��U@�,�R|>oX۝�����c:�c,�3��#�"����|������	�1w8AD��:	_�Դ���]���i܎[��ڸY��v���;���l�?�l�/T�  �ĶJM.����K;�a�K����!�û09��	cA �\s���xD�	ّ��o�.[�"���P w�������Ϙ�T��b��d^�-���d�g�5��3���{�.{'��$\��W=�K]J����yH~��gZ],8��Y�!�M��Z4��1�'(1@���m'[�A��N+4l����ƣJ�5v�KC|�x���[#Q3J��/�y�|��#�����)��bNd�!&cuK>c�t�S=QDy�����F4O��|��L%7�t��B{��̐�k��S��@M`yIM�5Tlo�-;�rc�ę	�f^ΟC.�S�P�FB^�l�O٩���R`��9!��<��z���r~ÛVqĴ|�9����$ �w)UPG�|p��j�YP�o�%E��{�:�G�
&�5��������Z��b?}��U��GS�u՚��+C��6ĸ,���{j��ȓ+@����� F�Z�I��}W�����-ּ^��Ct�����c<��x��&�Y, ��ҳ<��~-��\M� ���m� l���[���Au�l��ꐢxI�`bb�c6���v�јf���A��:k�['��{����X������mH���k!��ޛT�ӗ����~���yF���N`v[b�)��?S�Ό���k0�PEV�M��a�K9��ml���Z7Vl�DX|�/P�����~�g�P�Y��y:�H�2�
	�Ht�j;�J�d����n�Z1�S�n�ok�C>�@��G��Ţr`�?y�!  ������j"�;k��=���}P�:!ܚ>jf!���pf�o�ϻ-z�Z��C��B{~0m�l�6I���X	���U�J���2V�a��)���B���s�f��®�ĳ�6��� �r��;�����7=>�.np$X~�6d!/B�Z�~6O'ܭ��!��\��2�{yF�
Ⱥ������1V��]�U�	JBuBM��C�}kS"�j�ZB}�r�ظ��#�+q�f4~Y��ۺ�������:�&X�d߷n�����4��|�d���0X�@��n~`�˒�^_� Uu־�):�F�p�呎��iy�^��$8�';�%t;�he:��6h��8r+�*I�w��
����AWR�l�G��!t���@71\yh����Ί	 �M�c�N?�{:@��FYN�U��<���Õ��$��������	C����=�������c�*��`x����6�y��Zn��n��,-A<��_�bX������dX���}f4���m� Tn�x	�u6��E]yN�h8�C]JKp#`�8;t^+*���yxi4nH°F<U:X��F�]�t�hNڳ�$݌-4�/�x����Z �D.����?�����f-���t�o.u�G�^�e5���Ȁ� �Z��nn���3$������pD�'����:!."&e`��H�/���.��'˶����W��]�3���PE@�����۠�C���� ݮr�7p~��������l{P�Z�㘖���=m\+A�o?%��@�
�G�&�!�J;.�v ��`G����a7�;����Vy��J��,��oՊk\�����9�8?��@IH�6���#�K~N������8��GT�j�=5$n�hY5XzN3��i�یqȳ����)-��ق��G�/��6Հ�_A�bW���kOR���t�B7�Kr��_��	�zY�O_��͹6��#��cZ�#��휓�2z�ecD�/��-|�����g_��Ҧ���ܚ9�,L9�n�+5�&2�6)�̸q\��I��!q(�M.�$'3w��r���l��x���n��~9N���D�� 8���`����H���jx�����^�ƯM�E*/m��{�Z8H&�{��L;���I�.]�@/�z��d�}� dC�R�%��3��H�`���J�����-�X,�F��,y�;VqB<k6���{O~��U�!\�ˢ E* �J_r��9�<�VE�Ƒ͍w��3�zZ�!�B󅋉��8orS7���!��Y%��oH�0ޞ���g-g��������bȺ�o
�����D)��c����V����ysح/r�[���3vu��ć}�`�Eyh'u\��%ag���=S^W��*X�ýPL&6�yCA8+" /жq��/8�$f�)�Я�D�?o�	T��u`�!O1�P�飖�d˱X[����w��C��4��ݧ��qzЂ�z��8�z��k��9��#CE�S���H4E� \ʡ�f{��m���"_iJC�E��_P���%�*�:�I�Ơ�S!�J�ytqj>&�-ߟ�H���*��%�ĝ�F;�>�}�6T�z�I����4��^��j=�V�0��6�7#e�~v���}��'(�~�������H$��(����>��'����N�����`�o`󎒡V�I �w��mL�$B���A�5�%(�_3g�O��/\��貼=�jw�*������~����DfK��CӚ@5�>��&`�Rf7��)R�f�jr�fx�r: 3+FWkߟ-�6���	���]�ڸ�i��n�g��Mw.�o�Ǆ�*^ �v��.���]��w\ʳ��R���X��I��B���ړu2m�3Jx��_�����ڙV�
�q��un�l7��ٔ� �4i�p5�Cq����צ�����6�h��R���N�"����V(���XR޿��K�i��o$\��+�k��F�qَ��M��ݒ���_��k�V3o��	E�Z�����j2��O؀p�������򍩮��C&T�}[
�޿G�wn=T�S3-�Л��)6Kt*G�M?g"�;�r�\Q���气 `H��e>��O�H�"ꃗ�%m��!�+���GG�����GsJ��pК�+<rkZ���%-�
��Go�zJ�ɤ�m��h����ǐ���$���>�*�A�0F���Jl���?��:I[V,4�'q@�������F=�A�J�X}��}������~B�i�5�n����b<>Ѥ��ct
����z14�w+{�������+K��O�s���t��t� [6�o�,����%��H*[|yI�$�b	�	��Vbg�?z�4��M��ڴ���vu����'����=A��o�K��d�I1�1xjy�P�2�ќne�{1� ��w�`H��ٻ�N{	��M>�8�����������^7���h3+�i���<#p���3���\jH�m;w)=�L�[�Y��b@�3�BT�f��I@5�]fxpKp{��V]>1q
��E��B�G8#��&X����a��>��{y	Y�V�SE���-� U�Z�����z�����N�oY�����>Tɕ�뺙�x]�a���P�3ت�2@"����ْ�'�	��2�}�8����ln���B`�a?٨���˳FP���销�sP��b->�^�[��%��%A:'�S�����q���Ժj=N~9� �!�M�����) �݁b�^s����;09�;v��>�W^>QE:W*�FٜL�ߠqd�����g� � p�N�CVO�����/�7nV4���ާ%'����
�;�ľ7v�}3��KL����e'���U�u* z k�oĒ��g-�6҉͸�p�L�����h(5�2�����"�NJ��x�4B��[?R<F�v�W]+�p3�E�t��&63#U��2��s�~��`��:�MI�_��AT�4D���Q;R�B�U�b~���9D=�)�%�0���`Q���(�R�c����ĽH�����ŊIK �������������T���,�n����{�qc%x���bd�=��-S[r�e={#����;��Yn�`����a�5s� g�W����ٟ�ד��;VUald�m�ƕ�.�������q������0�Y�U��@*aO�FXO�V�����֙aaܮ�x�8>��﫻�:���Ww��sE6�
Ed�����;�����D(���Y)���Y�χ�o���p�)�(�bFov�Ob!���� _�ڂ����.������[�"���lmU�A�MNY��`��Q�BN�lR@Iݻ�?E;ChA���>?��9|6=�0������l��>Y��J}�tN�-�y�����3t��ji୿z�Z}x�{�$�V`�.���J��)8}"I��+J���u�qC]�N_5���V�m3��5��W�	�]�}�
���v�m�.p?�^FMP��bv7YLد	�:��~?���ΒO�Q�/���@�d�w��7���,$��|6yņ����/g5�������Y���Q^��8��<�S���Az��0D��U��3pM�֐AMʆ;�	�m��?�)a�5G��?��S�䍌�������+vf�8�h��9���y���-��ڎ_z�a�c�ٛn�A�h��EP��2^�PC#���IU�(.
ƨ��=[��[��&E$]]?��o�#��
ΐg	ZH6�΂�)�fT�!ڿ�e;�q�,U���1�Hz3��M�]d|V�v�f1n1a`?;�҂�C��qܫ��@��PDʕ��]��6��f׮���Zni�����)L����]W)��2 �h�Q��Q�]H&�N"��3!~�r��AF4?���`6Rx����g��#���K��Fֽ������	ޤ9-����'�X�X���s�����dⲝm���e�g�s�Iv���T�Hi�F�M߮��K.�1�3���pY��Av��/{!A��o���Fz��9i�]��>�X�x��o��M���KB��oڎ��#<�"�M�D������dHe����� G$>g$O�d�y�^[���v�h�7sͺ'X�UL�&�
� *��Ia=9�pw{: Hu��<B�Uڜk�8���w�O�fOG�t�;R�mHu��"3i^�@��v����y� x��Ժ)G#�j�g�y�'��PE��O�7�h�j�����)ظ��{�M��T^
�ά�a[9�Cˑ�wx���i�*�h	=�x�E-��cL�؀�]�z���r_�m��.�Ī�ŢVox�1�Zj��=��$�@���,�t6�|^@��[7��;hRTV�P����{9�
x2����pz�\Z���ٯ4͎�D���*nWJJ!���eC>_��?��c���}�O`�<�E��o_]A�[� ��AS_��ڴ�����F �aeʠ�t�5�nF�I
�8��V�f[i+/�[4!�����m��W���R��ɀ�"�`;ǼK���:�1�uFvj�j�R�A;��1?I�|w~�2����sra�gzy�ߩ��埈}.�P^�ǎ���5�#&x��	ci�Yz��u�N���k���t�^0�.1��;��_�O��vw����Kff��iI8�;��~+����=l���i������*��������A9�O1��]�$d�bl�C�m݆C���'I�U�2@�
�����#]�Kz��_��g�~Z�U'W��s�L�*P����B=���~�|HX��C��\>�ID����9��{.�Qs@�h�_�o��8����.hk� s�����V+���Cv��B�0����'����r;2w�I;1���1j�����k�Q�E�{kQH&��L��z�=����oۆ�] ���ȡ��C�ܫ՛ҷ�m����gc�cU���jg�:JJ �K> �W�7���D,B	�c>I�H��,��V'���=�Lw�*���c4�.4��s�~����]k�����y���P�vK-:�$���x����5&e�e|�͋�Ig�X�i#��3B�N���9�Gݚ?A{R���9�-���o�>6�b�MƖk�9���yk���7��8PSz���!<����Bj�&�v�np�76φ$E���"E<O���AP�˲?�o�F2_���H^X��P	.��4�`�c�`� o����c�.8����Ղ:h��|�y7x6��: 9]mZ]�i����6	Zu��Yi�ℇ/����Ӌ��B�GU�][X�f7�:O�M$�(+w���`u�>y(<H���
�i��!�[<�=�(~Q���@SM�����?Q3g/(W�vy�8�b��W�g鱍P�a� "�7DE*�8r;�د�����#��Cq�L T���|e ��B�k�5������Έ�MM���p�e0o�!mY��}]ō<D+�"Ak�EQ���<)�!�(SR�T�hhc��	���@�
�V�k����c��4�hݚ���wjm*{<ѿ�-��i`�  �)�c��.��̊���9F����S�Qr=κ����9�0�)�[�yP�Ls�`�@���Ո�.�Y��s!z�Q���[O��uZmH��Ӝ�,���tvA���w,��i;qh��^6�S�y�hB0{7Y�>d�@ۯ�%P5��O��<��Ŋ��\q���Z�@n+ w�]_�vM�؀J��lm�)#��m�^�tZj�#$A�[���&0��^0-郤�?.?�yI3�J�1�Zc��D��E��YS�G�dJ{ �f��ι��aG�C���nl�nAf����f��`�c���BK)�&n�Cο�f�z���|oY�G�@�ᭇ�x��\u/�����j��un��KA�~��s���b9-���(�~�N�j�r�]�R�{t,ϸ"{�* ��4��k!���I3Rǝ���V���1��n0��4��OQ�;�
�)�6� !�G����K�����}�t��s����7�^b�Ѳj��ثX���C�m����;ô��z-� �
��8��c_�PdVb��F $	sȁ��/�܍�:�&&vDԿ�?n�:�C��Ճۍ����o��ө^�QY&�W�jcL?��Ԃ�
�T�f���tM�ȶZCz�#Wp���ɓ���]�ː�;@����*P��gm�"�~E�X��Xk캎�;r��.����3�Ɋ�NE���Uu�uU��W	e�rc�@��Bt��3��+"7C��b�v��~�����䮃�R�P�+��?��Fm�Ah
Ե�UC'Ɠ��5��vV� �)n�SGWɱu�6����.�3�2-����d���]i9�ʫ2�^EC���1̟`Uj'�L_�
���Z3u���8/tف�@i�u&n?�26wJ�	�e�f8O�0�˺�DIꙑ��c(����'��g��	�-���IU�J�Đ3åX��+�q����~���'�RI�Hkl��]��~�;I/��\���S
������&�z���pDK�E ���<4̽��q��3��E��v�鷂�
�Y�2�/4�'lw<�s�)t�VK�_��-�
�s,��_����~O�^Ҩej���uX
"xem뫤ҩ�A���m�+��iO��j�i�����y�Kծ���vq�PA�Y���ڜo&^L�Xg�Ղg�H�ksА^Bw(uڥ�0�褢J~����&�����I�)�ؔ��ENlm�����(�R�&3��ys�R�4���^S)]Ps�X�?Q��P楄Y��$��M5� Z�+E�/Ύl��5@jl��n�&~:ʰč�����۩a���<���!�8�^�(_���s)W���H��]l�l-��Zp�<����or��<�ഏ�3����!���Oy�4��m�{p|t�n�k��U��n���eP(�Syr�O��T���B!��{g���~�R#(���>)�9~�HT�s��;''i�}�4䲽�^��	��t�(?���&�G�,gt���
��'�����B��sl���X_�WK�(�
���z&qi�er~��|D�����}A����RQ���&Rd��
�$��ak`h"����-U_�,�$v���#��O��'��A��.�P�u@p��d����I{��:�1cQ�WA��I���G-:Os2�:�]_ ����{���g��ɜusf z,Ek|���U-X��ƽ=
��
�Qӻ 1�uD��0=͚�m�e˟ݡ18�f�\�1*{�,aF�NT�[G�͗�%u+x?C
^z3�a�����bt� X �CU#�.��p��n���}���-ΜY1�a�����a�$Ɏ�
I�/U�S���b ��%�ݹH�ؐ�j�{K��N#�ft�ߟ!�;şx�1Gn�zT�X��H �og"���T2C�[�U����[G�0*�:��X���?��{��b7g6�XU��J� ���,A&����M�Wh&���
2:� r%�\!�9Pq`������:�ڂQ� JR����G���xSUY��JjpJ����t)Rޫ1jn_.UAAց� �-��@����@�&diDDet\������ ��T�I�Q?;�b�*��(�g:�Q����|��lC�bQ/A+�	� �ٗ����}�#�x�Y�)V)�;��o��3�X;�p>�ah�N=](jp� K�M�� �|�gq񸯿O`��3U;�(7��4��߱9ce���1���]4�D��l�F��8W�=�t�^�~:#�X�M��TTB[��l^�k�����켯$� }��Xm�����	�{��)jO[��?��o�{N��_]Z ��Ȓ"c����2��e���,�(:1���D�����҂9FX]��q�T(��+�1ˇ�ۨ��W�GY�n6�"v���9�m�W �8{�+�'��d�鶌]bo9B5k�C��$�?�lyRގ֋ �"2�X-�9�]��60�ިW�?�{�eRH��?�d;���b���X�aYIH�aA3����Q�_���(�쟦��TA6�����o�=��ڳ��F������."�z��aDYw6�
B���\U����q��M�j��W%,W��]sM�%f�+��+�.�������%������\�z0���	��9~ɭ���H��}Ё%^i��Y�b]'T��di!7A&O�CY��}cn60P�-]�K/Q�T�bQb�v���p8|���
R�����A��ִD�db�cO���7�G����4ݕmT7���^�Z	��)�)u���3�;���=�Yp��f�7��N3~�d����ͦ����T��a��}BK��E�9��в����n�w"��kpr6a�$AX�X�Ѥo�m�h��g���a���v�Z�йH����O]ЂJ��@���Ñ�z���=��+{gcPT��q[s��Ɖ�S7ʠt��셛���E6�'a����
�Es`Eo�8ʢ�p]�!+��:����_*�N�ڶ^�dE8���aV��)�:�-z`ґ��ڴ�?�>��N��k�3#l��5�惯!T�B(�9�(�t�A^�M9�ᾚ��R����ub�plPR�W�8�)8�߰Tv<�J �/h,	��V�|��ۀ�.��yǜ�{DLn5���Ō��\93�2�: �A?�06h��U�`F�Ζ!?�q�c����u����_r�w�(��[����"&���,�6��կ:���ZH�i�g�Sf�⋒)ߩط���F7�#^�ZT�[��=��7�6��������~�=#�!�M��NHʑ�i���z��܉i���g!���ú�B�,�/V�U�J� 0Bb�/NWҐ1��e#zo�Հ��Fr��LW+/�ȉQY�+>��y#�O��:ݘW�|�d���e�:חK���}At;NX cM���H`�6*�d>���T~����)H߮�k�۰w��)�M�l|�&lR�Z�.���?�7�b����œ2���m�gU���*��c3R�_�JAI�V)��W�V����PYM�W�e�|V~T�eٞ�'��^r�H�m����fsL�7y����#<֫���7�>��
�"K?�����8ޥܮ��6Er�A�c
q��zv��o;���΁��[%4�WBDud5�)����=k���;�[��F��o@�mo>C���/�����u�b��N$��ƎЯ��5���Fy���M�z0 �F�b'*D���C0�f/-^s�����Q� ���?�껊id�!N�Ǚ�P�S

��E�4��u����������h�I	�M<�hdn%Q�Ώ�A0jpx�R��w��/��,�⣭"�x���-I���}�$[���o��c�x�e��it��8�(��d9��Y���Eڧ`�5"���(��������`V��M.��=�:�ZYv-���>z�%>[K��Sw��~U��.-c���	0W����F:S�.�� X{�Mc�5�j�ih!\��	/>k��n���.|���*�ֻ�*�?�i@z�B��H�y���w�hʅ�y��D�9�Կ�v;��F��EI�����CzRn�v�BS���d	����m�rk�M�+h)��oo@�x����K���jb��B ��+�t��Lok'[%�vݯ�C��wg��%Pzc�o(���nY��z�h�H���z8�D]}��g��Ȋz�7~�A�6�qW�J�{��[1�$G-�[t�$�|B���d��f���L�*x-[K�lʈۆ{^�c�ߊP-��-h�Wbʑ}Яms[�������R��;�o	�3/RJ歷4��S�Iw�I&��`\�]�������#m�M�iu�^�P���Q��4p+a���T>L���eԅ�Z�c^���ϰ6���!��XW���;EJ����)���3d���.�����.��~F�!ѱ�+0G����Rg�{\��-�i4��Z�q�P�U��K@M�2;F����j)�ҹH�d��/������Fx�lA��7����u��@i������VB�Y��A#�����G����~���(�~A9f����+f��NwZ`|�|�ȹ�{�����b���~�te��Q�� �-�{ ʴ�)5�Ih����� ��[�
sG ��0�뱙�f�$�mR����g˯��#�a����|�>�qəc��|��i�L�&>�=K��4��z#����&	�^��'��JQ�)�<��Fj���f�%g���_L���;m^5�]��nw�������F��p�Vr"=�	,|��ן	��ժ�Ibo�& 7�M�V�˛+_��E�C"^1����~ N�S�"��ъ����#��O�÷sy�'�V%�8������Ⱥ�`;�*�	�4���խ�s��|��)8�ļ��!;����y�pI�?N���Ub��i2Lҵ��U$��1�-(�_<�x��η��z�Oy���6�m�u�����׸����`���:a��6�G�"����vV֊�8�X/wW����te��kܚS����-3?B��xQ���u5����H����3��/%�ۊU6ȁZǡ�"%˖&�H!�OeD��`�͖��o'��������,�(� �|���[1�p�'GΆ�&��6Q��L��$�����\�@�LR�\�_��^]�o�&�c�#���d�䠄sR�JE|B]��њ�y���[��(��P���T`bF\�����J�󴽠��r�H�s��WdO�Z�R�7J�N�OnN�e���m�$���3��^qޞ'�ԩ�'b���uep*��Y���/����������nL�7�4VLep����U��f��i�?m�0�
|���	TR�l
��"^��@-p^۶�Q�/���b&���e��߀��ڒ��������g�	�ex+L���T�4�����f���y� 2�o��h.]0��a[���{��c��}��$9߻��2�0�X��i���(�'�jeǣè�<�iBRư���-�g�!����*��e�r�i�JW�a^Z-���Ǫ����b�Y�wBV�X�c�XO�Q�H�Jt�$LC��DH0�m:��Y�@�7�i�ȋ�����Hb,V?%���)�I���p@%�|涏cM%��N��]Π"�dY\N��kD�:���ɵ8A�l���v��W'd,�|W5c�<V帇'&�m�I��I���qH��+�ak��G}G�1�sA������n�/�y:��2鿛��s�I��U�8W�%}��kB��w�/ #�Ѵ�����ϤF��vx+��*�&i�+ ���"S���x���o��f�)t���h�3Tĵ��H�ڒ�x+���� iN�7wC�^Lcnwx��VY%eL踜�k�)�@��	O�!D�.���u��N�s���\�����g.�Vr��Ugj��ZX3���
t�E�x=�������vH�w8����	0e�;&ؘܻHEw��.��e���s���˲��a�O�/�z8��=���Y{���Pц��ϳl�&��&�*W�����$��ū��ʅt�|=�{ﭤ뿅rV����*E{��b�W�N�Ȟ�D�u�����'��s�ﱉ��X���?�4Ζ��]L��=�����,?���J�R�obbE]�t�cǡ��&����8	�& A�B&jU�@-��9�C�I�'�t<
,ٰ�}"o<7�%V`��Pp�>>�K�9�.F,��q��!gF��I��{p�"��KC�t�?�O�h�Ҙ��G�����Hz3mi�Y@��=/C$����<t�@�nb���E�.��N���x���G����j�&��La�o+��C�=
�c�P>(ײa��,��n!`���n��t#|���Ċm���q#�ewrɇ]��J�l��^�j�WC�R�N�ݞ��U�U�K�R&7�J���N(:��ba*��1�@���;x5oA�:�vL�E��wm
��W������dx���r�W��n�6q�����)m�!��&g���-�kO�����S\#ܗ!`�׹���<m���.H�˃"�Q�x�do�&A1Ma��+K^Q^���e���-V�8��MrLPFM�����Q� =*Ϗ�?���.yW}���}s�?%��u�L��ˎ�����Vܥ �R�l�x|[�ѨT'f�F�j$d
��jf�uf��m��JM��{�6A%��|��0������wi������|ZU��C���$�)^�]�a�+����ӟ��WI_˱{�N�\�%%�&��8�IfY��̀.~~�M�������@T k���؅�@���-t-CD��1ˠsQR:��v;aq~� x�rƚIk�tԞ��l=��(�H��Ab.BA�sՊ�CR�^�x�u��Z$�&��[�ѿ�~H�����r��������$d�1(�R��@��W+|A�}-���J��P�U8����g4�}9d��#����C=k�2���0�W���@�(���FXtkU|(^��
MƔD^��� r�ˀ򟽠��̮n�L������2�ǀ���#^r�ݢ����ReG!ٞ�Q��żp̽��B�S=�~0)s����Y3��� �cf�8�U���@$ݍwj;z��P���,�\ m{�]M����(nV�^��Y����l峋Y��(O�/=��Bi[LL�Jj�籖\��#~��]��!�ѐ�Jͺ+%�l���f��1E�;��P9�FL����x�+�ޕ~T���.ʀ���:z�oh��%���k,��x���}���
�p�$��@�����H>D��7�l�w�;HD�j��c�aA�[	Jy�������Q��j�%5���V���|���:�.������OY�qY�SC�t�kc�*g���AǤ���2���Q���ez
A����3Ea����[Fx�X��W�9/$F��10�� �w9��%P@���&�t����
b�-zST�*wv͑��]�_�Þ�wPF�
��<��"��Z>��"V��?�2$�D��=�o�X��e�Yޗ3�U����օ��k�ā�
Y�=4�w��S�������f��͐��pAԤ�Eh�R1P�)6�n4�A"�b�`�33��E*�Qg�� �R}�U�&�T�1�n��q���5]���5�1�ym��z�y4b{i<l�q������Ņ �k+����e�X������Gq�balζ*����-�6��_�(�ǵF�F��TSXo{:s���6�7�z�X�M�fq��/3�>����6�-���s���J�R���e�0�ߠ�>��NUK!*v�Hs6_BAz#x�Z������]hN�x�����o�M���!�o(��y�f�|G�]��G�s��� �GJ��]6�4tz�!�5%���T���i��Hl4��V�����7}����6�y��c��P}�vc*���y��	�O7g��Z�T����t����zU4(�u�ymY�ʻ��J٧|�����$z�t�j(\�0R��j�� ����Օ�:s��i�*U=tPvF�w	�w�R��U�[7�����˄�Pw����Mzp�5�B}��pE�
�d%�:���{�G;�S����e�>o��@����m�|�2(yEs,�iL�A�?R�d][�v�r��s}�p̧K�\��2P%x�ז(�x�W lE�ORpSw��-U=���Ū)�g�_e�]����k{��L�<�0סJGX�>;���!Z@�	��V����M��X��	�\90;����-_n,Rs�3b��p4���:�q�Fώ���x�n/-��e����[Pk�Y��]龙c؇�s���Fҏ�dU���������fK'����!UC�����QH�\ܧ�3T�����ki�P�>���>�b%��dY��p
?��v�	:ظSX�󟑾g�.�����?t[�Mw�{�\z�_-�b�2ԑ���֥?�i�L�:�V6�KA���Q��辰G��C���?Q�~�<�>-q8Q�-��*�H�P�$y�̇f�cP�:�T��q���E�dh�mQ~J"�=L�����vb�aۧ�' Y�k�>r��'������X�0��vdTy�}��i�&T=[�ؐ)ϻ0
m�v��f�䜶\�c�Y�x�K��d���N��ൠ~V+l*n����h���w��s'�߬0��N���W����߼eTc��	"���3�g�Ū��9������S��f�iJ��g|$�8�~��ZY�]N�5Ȯ;�xf`�����O���/���l������-W�}�V��v6IsG�����Ujo茋î��Vݎ>�4���Tv<�ѫ�"�̘���uƺ�-����.��c�a8�M�$�芝S�,��Қ :85U����ڡ��$U�ʗ�0��)�!����Q8������]�����7uw8�L'��w�"ꦤ���ϫ�����4J��]ky� ]Ka���0�|z�0x-����}I{���=��?�T�����~7��﬊��ޒC_x��z��x��	�wŀ�-R�n�����})т�Ճ]�B����}NNjy^�5��X(�s�B@/�~���IvXq��:;U9�����l.�b�Y���="ʹm�����6hY�b��M�> �z���F2���#�:�]"��:�]�e1�ֶ�����$+�3#�o���3|9�DH�E-	��qy�K&!�E9N	�>��֚9愑.`j*�C��E� �p���q|9	�m�<�U�k0^A�aX�ŶTx�Ș��������X3�Ņ5���80Cˁz(����
o�=�G`�2'�fW/-�?��渡�3̒�G�ҒY|5A�T�����)�F�,��eܭ���i��2|l�2������Z��/P$c��c�b_CG.�_hiO�`Smf�A�����~]"�k��Xdxk��gdte���G	�Ɏ���=����'�ׅ�q?�1�o�*�/>^���W
�&��]���w��z^f������r׫O�֜����EZ-���_�Xo6����7�2�v�*$X��t?J�\�>g����ۿa�dH�I��ֽ .��i[I�d�}�l����t�O}E-�O�g%H ��a�>�\��d�K)�X����B���ۄ�S���k�6QF=N�^I������c�Z1Y�w���k�:���hY�sZ�[	��������|��)�A�i7B�
�0���ɛ�|�{so=��_*�h1�_f�hĮ�_®�Z$6́=�"�J�d�?Ǿ�4}����K<���,�dA��BE���+Un���Ŧ/��G:�iP�a�H����Z
��4 ��g��ϱ�Ą���b��W���)�AΕ�kZ��Ş9p>m��>x��	�_���),2a�I@��\X��{�)��6�v���#u1��HU��D�tx�ee_���F�Jt��ɝ9�y=PȟX-l�>v�#2,`>�4s~f�֫�ѹ�U�/e�A|P��\2b[��t7M��pT�%��`����n'�0^|sD���ߺ�x#]d�@�J$�<>>�X���T��22V�&�*4K���c���,�jh
��X���6�7 �xU���]��6�v+}���Ty��KU��9__����Wz�������rW�b)K��2�2���`����Ǹ�~Rq�#�3��j�Z0.��|�ߋe/�� �?���Zj'�'�/�cT�d�B%1��Sm�B�"ze�iʵ�;��뀱3i��B`�Pe����=^:��9��{�K�
⮖:`���gb�+fk�w���S��	];�ِ�T��tz#���b�r����Ř��ɬa�W�EO�ͷ�~鉁�t����(��Ga����m���oP��7۵�.7���(/(�lTӟ���M���I��9>�7�풬���Փ�`%�]�T:3E��43ޏe�Ib�2�a����Btu����ɧ��
�/Q��-�8/������\�l���.��#�-@���Ɏc���������?_��%�)��~�aee�5P��?	�%��3�����UW|=��e���d�$� R<��	� �8������%�N��&�$�.��\�EYy+�C#r݆��)�º�`FE�+���y�jfd��������W�����M`�jj̋=�F�W�/a1��5U,�-|tHHE���袚
�uB4w�E�*�%쉾?B+�h#;������$��>6��!P��'.[p�_h���A��%A!W���M�`�Z|
e����2�U�x�X���Ukλ{��.z]�$e�i����+$�P2pI:f_����}�k��<���L;i��U`\��&4��/�S���"z��P��ɜ�7�de"�|A�_�.�V٘�M�/e�6�*`�(��N%�I����t���+af���El�c :�]rِ���`7��=4��F+=��I)h��h|�L�΃��r����u���Iv!4R��9�{mxD��B���>��"4��#HU'6�e�T<AY�9��N�.��u�A*�`�$��H�~el� Ѷ��5ܶw%��X)��$��fY\���-Qq��\����<2+��i��l�J1w~�g_���:�)�LiW����:531*w�� Ux���ԏzb�`�0Yi9K���w������"-�f�B�������v8R���&5�<���2�7Q(�.Hڞ:%�T���~���Ӫ�ހi���.G�ޅ������!��Y��5RE@�������69{�����fˇ�r9��ֆ�G�O7�����x���z5)��E���H��a�-T�u!e->�b99����PO�o�Z�h��)iehp�Ł�"������@����O[h"70�c>�bIa�;�Y���WRxZ��l:ia�̪�� ~kڠ���4L�*�#�u�zE����x�#�L����ҥr8��o���&��ʐ�>��|��W�~�b�j�T�0��Fg��p��(:� M	IH+�")�C���(�����jo��DP�
��F�>�w���X�l��2�*������u����6�s��=UHS&^:p��z=��,x�-Z�u���	������lo��6�E��&��{��I����zu�A��/��5ѓ��w/e�N��8�2N��-�ᳮ�u��փG���*g��¯��?��2�x@Z��F`ʺy*e��J�6EJ��f���'N@�[�l�ٺ�d�Uf�^����f�ﱠ�%��2��v��\�z���Z|>P��b� �lr']o71�[D��^��FPl�����#Xs�혌1����{j�n$�`����J9༝F��8U�z Tª� 7px��0�X<Ό�C�0輮3!?]5�Ec��K$��D+]N�S�a�WJ�c�蠢�{Ȼn=�����2��@0��kNQO���i�:�D3�F3�-N�<�~? cW3q1����a���vhzX�	Ɯ��k�Q�1�:����X43��l(Yǭ2s�K;*/j�pJ�t@�	�ymvi["Rg��3��xԽ?uS�"'�R���x�Q����(�Q}ՙ��c%�|��pB�ϠJS|�|�h't!~25O�����^�aH#>C' �����@������VVI�
���x�t��q��zx�φ0�'A��w 2��|�V�S$}*V]�y<l�����df.�_�	ʣ/�PFYD�z�?n����KЬ�Q��>H�˃8Ʊ�g�Z�7�z��!�㖇�m�s��;��
cߨ;�K�t�$@��5���{��-RE�ZZ�?[GG���|���D���@�,���3�):���g8���X���`.��~�L������%��m{��:��
��eT��(,:�:�A������p����"�$���9�s(�V%8u�:@��e���h��R�q$��5�B]v�FM�R����k��>�S�s�m��)*�t���*u^p�������ǟ�"yl��̜�@���f��
j>IE�r3�7�G��DT`��D�E��{���� ��ħ�;����j��}���)e�;���Z4V Y�)47��mܮ�|�߳a�6�
uFm���g/Ň�Z�=���"E��'#�����̅P���W6J}����q�9���KH�@]�/G�Q1�w2�@�	?a������z]���Ru�t���;��g���T�bg�e��D� �<���[$}֬���n[�LG��iX"\n��S�b��W+!�䵖�r�:�[+�me�����mVy+�s���Vqx��י��L��B��3g��":>��ڳ;��U�T�lp�}h1�*�
�2hI������5���� I} �
y%m�Hޝ���M�n_���bNT˶	.ok�
j����,
Ϯm+�#X�P�����p���ā~4Yi�$QN3�Eq*o������r�H�~B�J�,�����yH�'�[f����#��qqpԻV�%?��W�J !xf������0�����0�b�S\J,@��u��2�x�zcv�zs�쮺n�0�Mh��,.-�O���r�Q�h�����*^����� ��7�gI��JG.�SK���uYm�`�5��g��4���h�:yZ#�c��,_� D����#9��k찿\�F����X�&�
�����~G-'"
�픸5��g?�Q�����<^Յh'�v1z�i�pV������o$�;jm<�p���ei,�Dr��v2�M�l�zQՀx(���h�-�m����:%�r⩟����7�0��m�>�5� �FZ,�&?�/Q�dʕ����@Cm
i�+��v��ځ����j��D(���Z0�j���M��h�1E`1`0{-��.����I�p���X�i\''�nn=���H.]��ʢbz� ��ZѸ
Me��!�=��Ōb�����F��is�-kN	��ɏ�ļ|��pwh�� ��C��X�C����y.x�C�HP&*	bdY��;��!���qn7Q�ك$Ϸ���M���1R#��%��N����j�g���R�H�f$(�b�\hl�a=	G��Q�*�
�)5w休�̙�'l�w�m�j(�G㶐��2���2�^�V*v�'�igL�:b
��?$�i`�?���!md$�i�Y4BN�(	��zХ$<�-�RO|�*�|\��t�F�Aa8R8]�"wұ��Z h�[Vye�e׶0�_��6�*n�S���&3U��0�l m��lfE���Xg�MLp��'����N��-x��*�\��D���W������&�E ����W��b>No5�;���=�!��n�P�Ш&0�0X/�Y[cM�@��?�]nB��
�v��xM�y�e*��s?Ck	(k_i�Wj N$-֌[�|h�>�z�6�W
3�@ ���w'�d{Yg�a���q���xD(-z���L���ڗ�%�F�,�π�m=ܘ�[}��sõ5���@G%?��P�jWx��[jƈy�Ɏl���R�C��@l�@�Y�{V�&#'
jx���n��=�[[����~���b��]�!��`�֌+�����O�����5�T�͈G���@������܎�-L:���h�`0�������	��*���L���4��ջF-p�g�"(�[��ԕ���"�����Ps��y���L'HF�M�묞 �ۡcfqH�pۯ��F	VB��AV�̦?mp��"���M!�D2��Sl����(�gp�&���� �Jܥ]��7y�c�>��O��P���O��$>�[��ЛЌP����\��k�J��6�ˏ�>��|%�P7�W4{� ђ���7��)�� 2~G��r�?���+Ϥm�Pjp�,�Ht�a{�;�7sa�lwC�g��c���$�������P���SAf���D�	���X�zim�2n�k��5!�a��dzՈ�%�B�yڞ����1��}a���5i'��M�kB�M���V�;3�h1�ɩ�"yef���j���_n^{%]���h9��s��\¤����_�k�wM�D�K��M4�F���_|+U �ʈ����|��c�j�?�ԯƐeUs�k�K#IgXD�
{�<P֧�Ix�LP�m��
�Șη�5�.�k����s�����s���}޼�+΋��f%��73��l��l�ʶ0w�	v�q�t��� a۲�1k&�OP ʘ{���}�Ӄ�u.S�'��@hM5F<�������L��-���h�*N�`t�9Wg��i���c��}N�I�{�m���62M�����f�\,�)�x.t����D�.�k�߆#���K�Eo��JP�����"Y+2Z"R#��[-8�^9[���ֵ"r
���`��,�@����?�$bEc�z�wO��b&-S��)�֊�ݢ7���kֆ��f/T��*O�:�S���8A�p��a��5��X��
�6���Q�O�^�47K�T�y��'���}iK�ԁb�G�f��20}E	reȃ�Xua�z����[;�$�Ր1%z%0�@3H�+��6nAb��0)2����D$����aĻ��/
�}��j����۞�7���z���M���\U�,���*+�Ѕ��k�ʇPo�8��Z_bKN�L�oUr�yΉV\�y������T���c�t�-Vv����Xထ�s>\ϐk;~[�G�b3*^��0��5�ǎ" ��C=�֬ik��p1AlBR���I~9v�R��#�9<�P�ҥFIW�'<��n��Oy��k��a�(X[Y��m��[�����ɈK�l����1��-2Q^�!����Z��*�$v=v�#wӚiM�"c*&��";�:�m������E:�EA��t�ǁn���f��7)�!vl{.b�k��b�B�<��w=��@���z���>^#_����(ʆz�Ņq�fW������!{��t�VO^� >m�b2�c	�ӌ�(��&�ڹ�R�9aX6^i��掁�]l���A�-u�sE��&2�R���33���~M����\Cc
�����S��P\�b��H?���n���*!��=�%��(��xgu�l�?���	���q�]�xy�ǂ̥/�m+ի,ń�#�A�i'g��G2خ.i��c���#+�S,�}-Y j��` ϕ��N��� �)4�BLޒ�Y9�$pi�oY�dR�q|�fq����?]�8Z��o	���@)��-̧�/�h�n��|�g�HjZ��ٌ�y<���a=/Q�aL�GSS\D�]�jE(��ķ�m-l�w��Z$���~�a>A̿��mt�)����wp��0$�Y��C��@{��d~��y���ż�����#��N�n԰N_i��9��)/���nd9����E|���*�2��i͢@ñ*�kz�ѓ�r����.��"99�0�Jf)�a}��GpW9�`l��6-Wml��=��[�;���Ý�ȕ`��O�O���ћ���L�`e�����D#���_���4�\�6ۺԭyY�8����)�_!|�m`G���h9ӹ%I������P����Q(t������]��?��R8l�KEi\X�p.�T���@Q�P�%dy�E-�4��P��Ɛ��9S)!�Bt%e�^7���2����
�D+J����%"��]3�FoeKM����:(����c�l�$���'`���t"� m����u�c�*�̥���)^To81����a�bX�� �����j���#v� ����",o`�1:�"R8ƾ'|Qx+u������.�$.��"a+��3�Q�}&�Hx��P�*k*������[�h]�������B!�Jz[i��mu���S�雀т�R����[���i�����+��*�=>c�����3����b��<��O�s]�ɘW/��|�Y��&��~�$�w������%i=p��7�֜� ��
e�'P�%�- �+(l+�1$A_��Ae�O�AA(�3�.� �1r� �F*�R���
��"�JKl���O�}���SC]'m�2�c���� ��l~�H��,����^ѯ���QsUN�x\VD]w������P|�RZ:gD8U�;�0��骰	R�Ϯԫ�qϐ��
4��Uc��3���^k�cp����m���}�9P<���������? �����BX%�	8��i`i�`�ցē�Ki�V�������л��M��J�U�t�e���C���Ҩ�P�Q����*8�R"jB&`�W����}�<��e��n�A���'��c�%�fЍH�ăP�CZ���^�E��΂�K��'��� ��m �|�>���?L�@�if1�����V�k\a�~kVh���A �6�J�� ��7T�_�����2�U�oY���Y�k:�Q���&���˭B�=� iY�h�5v�E4��j�,�޶�Z���Yv��!��9�]���F�]R��g���3�mF��׵l�m9��zS�Zd��su�xEij��*��؉�R�M�Z�-2E�<�U��i��)r��L��R�t�ݵ���c;��o�P� �d^ٔV(�9���?Q�,�{K����&�iJ�Oi�~�5,�0��轍+�~��J��
����YzZGbK0�ղ88�LjG����߭|�|�@2�!���ps�Q�۠�C��.�l��<`rV�� �`��?��7$lk��:*�x9��B�7�َwo������"�Nl��Ey���o@���Ol����5�H�us$�B˨�Ǫ�N�'�v^�zm�m0�Skmj?�J���jW�c���z\�Y�*4�\���Ǉp����bxAw�]A(�ݿ�r�4��%��{ؤ�-�\ʙ�'��Ŋ��]�Y
�ꂆ��t�����R!�>�u0�
΂�펏):���}R�m~]��E�P�t�<v���#��U�w�Y�A_,�x<'�&�K��0���>��0�Ƒ�T/	xke��q�1w�ߠ�k{��P������0#Ĕ��gL4jv�+�s��f�4d�=�v��N����Am�Rf��;��Ѷ�&Ȼ@�Wg�@w�����i��hHƀ�~�P��sBY�]�VZ]�g^���L��[:�������������с��M� �ym�zvrć<��������|x��ĀS魳N'`,��>�Z�w�������f�����^�rp�YIV{g:0���'�CÇ����8�	� E���'#O�\�d34L�k<�-<oo_�a��X��2����@��o���y�8����(����A�-���ö�`#|��`/�}K��{wN`��]{S$Kg|Ⳇ�vB���eE|Pb���!B��zq��@������fв�-/G;!��Yy�` �CN0R�p�"�R�n�ޖ�����?;3����{=?]h9|��Q����Q�Xx�U�B���/0_�Jw���{
V� $̢�u����h��!�����: +ez=O�9��߹���k����Բ;��W��K����!�i����Y�3�A��(@��������c"o�yq{F�r?w�g�A��e�`��-��pn�z�^k(1�zI�M<o�$�~��������.p^w���$�v`��Nû6��r��^+!ڹ���n�<wC,��ђ���uaI�x)<'u0���L0&�m�����W�Y�M�Gl9�ϷAlb�ָ|�2��ʹT:WI������Ӯ��������L�i����\ܚ>�4���C���A>��$�
�r�z���P/[>BV�t; we�"�A���
4��c�.��(��z���{���� ��bv ��*F�����jԻ�*�;b����Ks�%���:�؝��YPtiW��g&\D��_2�K`�i'��c{x� 1�6�q��*!��Ҫ���mKgU������'_��(-��Q�Te��CAG�q-G-�d������ͣ����j����[Lf�G�C��H���zX� �S>`{(�J�� �W��i�����D2wp�
��"���M�n���R\�pD>j5N��8��˖���0�^u,<J��N�N!^N���$/R�������*�Tǖ�S��+\׳m�rjx�Q��:`K-a��e��"�K��ɟ��2�B%9ۇ�v�<q�W)_�2�§��	0OsO����x���/��	&2l�(N���W`��	fU*�a5D<'�u��$�R�!���ƖZf1^X�p읩��sD[�WB��Aݩ�.2`:��Κ4�"���Upӹ�ɍ*(>z޶d +JN�Lb�(��%gFi���5�F�m��j���#.��=��	��:���̓��$�������۩k�_~�6ߓ/A�-�W α�H � F�&��t�\<�^ �"�
�Q���.'��J���\�YkN�ư�PIӞ1��Nh�!���T��'�;/���V��g��خ0�׹������|M���de����8�gB�/��"����ds�H �j)��d)����Y������(<s�$�cNE*^|q�11���$��܌ꑝ��ˁ,��;��";
z��Q�Rl�ϝ"+[����fMdߙ��7�A���kO� Uc�!���	.&���DB�$(��m�u�{H��XA`�}{{��:��e|H�^.�f�s�)�Z'�1V�x~���ת���z(~�ٷ%�e4�OA0��V��D�Q��$����i[B�/�/D�(�� K#��_��l�J<�D�.u;�h�;��x�$"�?�#�=E�e����-h�CTvW��f��0��*�����U�*�vR�K�&���"yv�!�}ݥ�\_��c,S����}a���-��4������.�F,<��? `g��[)�|��g��u���5�͋�S��&~�Fo焳�gAj��E@�+��`$�P[�t)`�Dr�laEp^eWȵ��R# d��h �p��\d�@c-[w��tD�ȧ}|Qw��[n�K�^�/��<�O��n���k�&�v�~E�S:	�`OH���s ���PD��-+����� F�vF�����)>�:�JM��[au2�������m�/r��c�!���)�An�,�����pv�Y��Nݙ�@���[���ҺgE�����l�h��q{|��j�ױW��Of��W}���YN�ӊ����k0EZ��)/�!��#�E(���(��#y��V*g���]��Z�NY!d���N|z�h�f+��]ҙ��-?�Cދ�y&�B��vBWg�8y~ `v���^E�܊V�y"��=~j���^�~�Q�Bj��r������zU���� -c�0����q���\j,��B�Y�n@$h,���#��nnZ<迓2�D`��$ .�,!`�&�g��.�HuѼ�T�6���"�'mnӎ�ڠ��iB9�R�T\m+��205BK�A���_	y��I40�б�.Qʼ\��n)0t��jٚ� ���,����~~�lK���T�l�떶n�53_�{��n��"����5!�UX/#��xQ�W�V�,�b53��o���iV�:�c�`ji�m�~�F"s~�^�n���jِ��Pd�To;�q�_�'�A�c����cz�~S��Vy��'���=�]�9!NTd����� ���˜0@�"�e��E��7�o��q�H-�����6C�$��h%9��.P�>�-�y#�rC+!�a�9&1+l�l�m��~w�=.|6*h�u{*��oG��j��.Z��R<��cF�z|��n�g�0�����������}w_��)� �p��ae�C3B�*���M�P!�>}M�+%��Մ\�gaױ��Ȭ$ۢ�+���������=�:�� ���$�\CE���G���H��ޤDI�tD{ŉ�0��B�$�$��JQ��(��ΟmŰo�:�Z�R�:�%=/���H�WP�_(n�L���Fm�U8� \��f�ǃ��Ӵ�����j��} %ۏRrm��}ʾa�H.�%��CLBg�q�9�dM���La�v�4�Im��+�5�����#��`�����w6qX��p$�ǪP�k�����-Z��,���ENB��AlYJ�b��Rr���>��c12���P ��΃w��9B�	���?U�2�p&��c狴�pj���l+i��K���ˢ���r��D�7��X��V��T�5&u�Y�Ư�Y�?m#?��
C�P�}���ˤ�3��p�X-�#�A�hy�C=#k@/]�"ҷ�	�������_��P�FB��W�@'��0uA���ױ0	{�wk^7�wz�*r\���P�f�.����o�,l6(kv��.0qlu���2������ �<5؇�^�k �B���mk���2X�&Ĕa��4�+=Eƣ� �5z��΀�.��qԵ�}��O��
@J.,K!)������p7f"A��6�0�	D�Yw�P���Z�! 8�z^��"ڠ�?�Ao��6\��h�b��s@ ����\���Y�ror��F�U���>7!��*�t�f�Jkֿ�uA︔���<����M���'ڦb��"$����c50Q�Hc%�c�覆�����茐,�4ȝj�i�=o���Ȃ�=o�ڵb �E\g�1�/�A�;##pd#8,J�=�}δ!��BI(vQf����G��DO/�m|u�/�������޶������gi����%��Z�d`�|�tD������)��w�8�E�"�Yޕ�B5�΄�f7��1ά��TL��t����NB�-����Q�(��Ɍ��6돝r]zPC�a�u�1�O<_ �� 5�Ȯ��C�ض;K/�9C��n~͸n��z�mx��,��g`p/=��x�0k�_��ȳ+�n�B�8������p ����]?MҞiA\���)N�6Н�UcW&�/���`퉁��)���D�e:�^�h�\���<F���e��?�q;�I��;Q),o��c�RW��?�e$�߼�<R-�� ;re��b?�z��kF/���ֲS�ݎ�8�σ�]+a}]Z~.�)+llU�%"�9�1����ᄈ|n��l��&���$� ���3�:�������,5�cM�!�v��?Pi:X�X��
���Xh��t�$��E��� T������Q��i� ���2�1����&�\�^^��P��r8���������Z�<HEF�Ձa��A2,�j�2zJ���u����&Rm`*��)Q��p��6ɗy��}�8���E��̀fo����X�wmyuL�<���"-~�R�D[ev�ͶS=�kN���������jb��_D�����-"d	1'��5��B[��?��wF=����C�AqT��?/��>|Q�d7�H��+q[�hVF6�X"�.��na�e�����*_�Kh��J���R�A���Q"N��\����Z�1�.P�r����������/�����#=��Y�p�F]�=rɑ6}<:����I��H��OCv�윳h�@����|ӶL�G��_�1�4�5��$Г�_Z&5�k��}�1�EknZ��|�&�=��Q&�~&#᎐y�M�UӒ���x���oi�|���eWԬ)�|3�*����!�a ܼjh0��j�@;�M:�pn�����^}������{�A��O<'T��Q7��I�F�����'���;���<"Mb���63�b[&K1|�e!�0f����0�]҆՞F0N�A��S�������2����-<f������B�%�$��q(�컵x�S��ǀ�-V�A/�E�O��28�-�U"�]�P�t��n'D�"����5�/N�ݛVY�ڢԈL�RO���� )C�1�R}:�ô�R/��v��ܕw�9��$-Џ��\�A��E��=�TܙK%0�d`�����Υ����#��/����� �W�%f�mK�1PHj�7T�#e.�B_Kg�"��1b�-����l�
�<��hn�Ц�w
���a
�^d���ʾ�ə�L��o�4�޵���$Fl����/�����@oBԕA7�C��-:!e�}��<�j�[A���%'p��Fcy.��-T��I_)2��u��aG��(׏"��r��#"��Gز#�s�w&�|�O��RY������E#��v����*vۛ��v�~(*ˈv|S�tG�G��K9��t3ߋ���>��}|J�o7���|ѽ!�;�*_�A̼W�h���?mE-}��\G9�D���^����H(SOWJ�m�Sl5��gcڨ1�%ֽ��Џ���գ���S�.�jj����B1�>��j����Z�14�~��+h'/���������x[ru�D���`Z������2Ly'[���p�b^�ʊ�_�mEȻ�s��}��l�s�:�l� {N2[�=����6_���9�_\V�H��I����o�sz)���3=��)���\�ᣥo������v��$��2,�A�<l�t�[��'j�a���Q��}��L��=~>I��Xk����7$% ��{����Q��t(�x�C5����.C�+d~����.�kI,7y�|����U�����31��v���
��?	J|�+5���0�QTvY�O����IM���z�����kt���T��K�tۅe�K�+<	�Pk�ڼ���.Z���#�v��:��ܺ(������kS�U40�[�#g��QCx�&MtV^JuB x}��p�|%���ԓ�1�|_��A���^:��OȤc'��\�����AIa*�mtV���U+*z�����Y�p�AM�H��T>q�~8\�Q�佃9`w�l��[M�XM�e�i�c�����h��kâG�c��+�9mk%���+���;�aC�
�UY_���4n� ��gF���U(���A���v�@ݜ����}��"�6�)F���E���v����	a�Ss�<>�Cq#L� �A��FhQ hKƠZ(���p�1�j��)��a�W�q�xq�a�)���2 ��Z�z���J��N5�r�sW��,RìJv����ؗ�x �i*��(�������%��`B��ǻ^	��2��V)��K��	�̭��+0}��w�ų7#��9Qg/"��Bu�r�ݻ؍�u"��7,� B�?�U�G�MՇ=��ٓ��Mx�/����'ꆔ�?-[f�߾��?cIހo@xE�}����_�]�~"7�ks���VM#M]z1��y�M�Ft9oDߓ~��Y�SfT��w��6�����D�S�[Lr]]�a$����R���Hg��9E����U�D��f� �Op-�	8r�Up*�p��8!��8�Zt�P���U�}I�Ķ�3@��-]�(�:*B�?zrG����P�Azt��j��jiI�ԗ��Bt��1�s�IU;������5���0�`!�/
¦��ZՖr��>Kd��maZ���Җ��|�4u��7e�:���H#W��!9C=�X̣vxk�ǫ�4V�_X\%C�O<�f&*,r�<t����#�t���P�1(�-�s�a�Ma��H�;?�qS�i+�˸}��ھ��D"��ˉX�������X�?2�.��Fe7^W�?�Z2��O��'��x)rT��ӄ�gv��ګm�9���Rºĵs)B�,��&�	\9�F�s�
��/�R�݆n��tC���r�?�\S�hv�����S@�v�:ͦ�A��˭d���4M6YO\�H`��$��S�����5�����*w���W~5
�@�)v��Rj��c�I�>�[K!V؉��wޘ�� ?��V��f�Q�:�L,^7�"����F���S�t���z�V<	��Üo6�Q�%ɧ뇍��!�e���>�)�"�5��}���<R,zJgE��l[�ä������2+��Q�FA���AB�q�c:L�Z#�8v��l�M��G�?M�aE9>YL��?5���(�W�K�vIn�-ҕ!��K���-1�Z�tuIz��K�W�*�������y��ϼ�+ߢ�.Z���& J�R�/v0U�+D%nkTr"[�(���#�9���ONo�I=Qj�k��f�Җ#{@M�����k^C�e#��D�����5�e�k��
8�w�.䶓d��n��8����Й��j��?��+��,���Ȑ������ω�2k�5��(��Ӹ(8�~����o9`:b2����Atɒ����b�T������J�����5P ��[S_�Z�Ĥ1L�����z���+�� e����]I�!>��a���T���|�K[�Mwh$")gz��N�w�Z`��̜�Cƹ�o�Dq%�z�����N@��P��	{�	K4;S�z�6��m��q�vt�v��v/Vp���lrM����3�W�4�)_Ж��}"�z���LR?`m,��� I+�Pz��̂�K~�x=�x�ٕ�^F˘ZŇ�A�K�q�%��H����y��{nփ	ь~�ң��E�� ���u�ɻ�$�~�Omq%;�#�W|�H�L�S�6}A���Ġ����x��<�	Lo�He=&/2�g�+�dBs���*��v�B@��L�q��Τ��_-�T#8̍��[��nj`���ӳ4dS�I����w4|3�j�mϋ?�]�/�}�g~n����5.�;~$ ��:��	��3�ġ�D�kE |G��k��o��s�N��XA�?��?,��R�4����jQ��{�}5��;n���[�zsX��Q�xf��ʳ�U"�҄�n��=<SR:m@�.��6+p�GKv�]S���=��T�~Uh�f�9��۲s�b�h�^��L"��2����W��,�<�g�[����%��4� ���[��ԭ��;t6 ��8��UY}L8��\U3�������p�֎��傦�S�V�/PSI3������Ç;:�r�4_t��F�V��U��:K�9&�@�QC���,���>~���=�wQ�߉�/v�`����0a�Gs��5��C��eZ�1|#�AQ�-*�b�%h�?_��
�I���[O��\�Aj>����.��WVP��JJ/1B"��#����0{��'��,�=33;�(�^���[d�ȼ���^�DJ��:L����6�O`�ƒoL�Kjx3=�?&:[1J�k��&3��6��� ��
�ԫ��4�*P���^���c\�w��,'����70P�R�J�]������TLnٞd��'���ܛ7�^��<�,�s�teĭag���A5>Qm�Q}��+���G(*�S�Ht�-�6a<��
����9n즁|�y�:۟c�`#�&]��_!�'"M��6�%q�ib����o1�E���kw ��.�Sh3N���q>B�ol����gl�#0q�E���=~�zJd�uO&+.KfǓK9�R��َF9�hĽP��ij?�>V�
"�Q�:��}��U���ڵ]���������z�$�-~��e3˯�
���˟"_��L���Oa��Qk�kz.ޠ��[�n��x�5��W���d%�D��K I�A���5��e���/�;6l��+j�[�)܏��
z5�wӓ��h5&�%7��Zؔf����{��#�$i�}~�剶�`� m�~��v�)�>�?g�U�0D�\��iHY��68b�:T�V�x�"�o��ɘPGo�>��$"W���D�1V\O�����b�6g6�����nF��R�5}#��O�M�>*��D��h���-ѡb���F{o�^&VoYփ�K���u>�0.���kT��+Mh�+�o��/��G���Xif���/<�v/��s)�䊜����a� ��f� �S��!����(a9Y��^��Ի���4����v��#���t,Iu��A��ɤH�=�ѡNG���c��Qъ��('�6��P����Xn9,8�/U A}�V����}��:JlnGW3F���^�8�rTN��O(ҩH���3)��q�:ݝQ'޵��Q������p՟�R��>u�
���jKX��Mj -` k#ݙ����C���"�ݵgu�!�5���f+��X2�%�aI�W�'��A�)��G[@��ʉN�=h�}����8�Ղ"&�gW9/J'[ܩh�.��y=�L~��P��7ōL���������v��<���w+ dfˉ�k����J��@�i��S��`�E�=g�p!>��4��uf`�.���Nd�	j��Ԗ�H�f�(����O��l��V���ʽ��c%��MS1N]�R�.�AA��k�����!E�ֿ`đ&���S�	3M	�艤������X�yF��5�8��n�~��.{���+Q��w�ۻcO����q�1����یFߦ����(�0S��?�k?�1�ӨN�}�Tt��ҏ0C}�����o�A���M�I�B����<��&�����m�c��!�3�j�ۜ������@G��4�V-my�� ��ʉ
3�Yќ�Y�z�4Z�d�Nܛ��� Y	M,�.��I����������V[��Vl%Ҥ
�ֺ�j���8�����w����u@{��Bg*�RY���}:a{�$�
	�(e����88]�9�jX��'~{%z�(
_�1�8õ��:�90�B��0JG�@�B�����Q҇/�-��f�O�%>�X\נ8��
�W�W��2���Zj�V�
�o�`�/o\��s�Lޥ�j�
�ʑ��z�h�������Ɯ?�f�U*��o���[��eha���\�_q����L7��m:N���}]H�h�k�������8v�rclP�̮�Q��{O0.e���S.�RNց$O�����[1��E���b5�Yn��oUF��r6v�1��5}e�,	��� bN�{xF~)�� ����^( dn�* ����)��1��i�?mo�9�����cg�Zy�$�6V�:y]�	�P�'��ʐ�$g	�`�eˉ,�(�p��w�I!+���E:�>�6̫FG�x��k�6��D��~�@g�u�zJ��s�쬋V���q���J�J�E 
u�#]���y�`ዣ�	T�A X��t╔�D@���#$.z��4$Hf�ӟ���g��d0U��O��7�t��*}��I;<,��!��.�t��e��w�AIf�O4Rܒ�!DL6~r"yEVY�B=ڵ�Ɨ眃�o�P����/#e�.��B=�1,�"0ZÑ8�|�LZvF>��z�*÷6.��u2�?髍H��	o��xE�Qf�[a�C��
Ϳ��K���T�Ȭr�ȉ��h떐�� &�A��p�����ǌ�35��t�����'`Rsީ�1��A|U�}4F/��L�-.2?1��6�tܛ�n��By�V>���rmj�C_n�W�Fo���0+S=e7�x���hS�R@Od��D;�1U��*�`��j����F�'ݫ�k.��G���nm�3g��A�*>tj�h��c����$Y���[�P<�|��FFJ�F�q�4�a��V@��i7)WGW>/b���X��+e�?��xV�~žr�Y�r'�O+S�H��۔���kHG�v�^+���:�&:�ھ��%���fI?��!!nu�����������Bou�f�rN�<+4��hfy���7��1�у��R��j�� �%1��}�&I-r��*��I�T5�C��y��v������E1���c��}RS�d��;!�s���8]�d��*˚9�]f��"�lx�R�=���U��ꯞ�\�Ѕ�B#L;��Xb�앸�y�7��v���}�0a�`��9{y�÷X����õ,3��¡Y���^���(N3�	&��c%:>"� �bcN܋�Sd��ujh|F�[����2i��ry�&}юuDh'������yQԭ�q��|3�q%:n��8T'<���F
%�U7v�?� 7�7���K����*cVO+��*�	͕��B��>w@�<��PG�S��̎�"_I�E�����L�����	 ��K=���Q��L؟7�G���
�B��� ��Tdc Y�S�G��׶Xl	˧�S�l\,X6�����]���l�t�T���R%�4���Zj���s7�٥��ƪi�I�ޖ�-Z$u/x���9(��
���[ѽ�k¹A���DUh��f�.���Y��g��w���]N�NK��w�﷧J+��Yڢ'
T4�v@#��%������Uq�^����9B���xTU��Ҍ@ߨ��S
	R�)� @lX���[	7�	���O(Fh/�j{ٲ�a	�7vm�]��N�[vd����M��߄��lM�;'G�[���qݫP%�(kv��	��ߨ2Ud�
vψ�2�
Fi�����Ra���g�&�0�+ع<�Y�|�����`K;Kb���Eݴ�</���*
-�%�}˛������/m�©d^	��w\�d�IU%�1��e54;����T�R2�4�;5w��x�k���5!I��3t.�C������q%��j���d�˚�]�������Ƒi�� ��.��.��<u(�)���^����5�KNvS�碅��g��!���>&��9I��L$�Z���߀�!����9 ����
]��OfM ����\w?
�����?G�%xck�1��s��a�Y�y5f"���V�40�m����}���̻f��O��?�Ι����(.����=���~�­�H�-�k�+�>0��(�L�l�쀎���`]���ek���$�]Ƃ.�ҖS���o���nSP�E84D�ȹ�榮`~V�p#k�~�B[="J�)!O�<�v��ҩx*�IໄJP��y�o�C;����ݴ�c��}����d�6���0;�C㾊���j���b1�o�S�>�K���1큗n�j����2Z�l&�v�O!�iTD��Iǀ��y�G�A��O�\���dc̞�ܿ�iR�̮�*璏i}���y�\	�E�k���Ģi֏"o/��F]��^�s^��$��=�/+�K�4Lt���I�O��(?��[�r����DP]����b�9s�¡~���1�\�hoH���_7 !�������}�E�i�:uO��
�Ra֐��HC�z�IR�N`�셣;�O��.%G���f����"��6�C�"嫲�>HE�i�z��j�-b�:@����u��ӻ�W�; �s��hu �r�qm�g|\���s ^�=�ҷ��b񇪤���~a<#Ū���7����.�U� :�6+�3�2w|竼���
:���J��H�=��ѣN$;R��N�i:�A�7Z��>F�q�!��SV{3��<&��a/>GyC(�M�9��O���˨��c,�dH���u�5)Lڙ�O`�Y��+�$�K6i_�R�,;n?��]��c�3�1=FQa:�|��x��&.�(�,_��F)������s	���
B�����������[��
 `���sq*�u2�?�e��P�,[����y4bw�d��_��4I�w�@HD��]��i�z�i��q����O"��.\���VR�`~��y
s�$c�ϖ�C`�R.܊��x���T#r�yP���J��y�U�I#,��z�>�q5NY��d��Fʎ�k��g� {ϔ�w�_M�La��?c�]f`,��A��Ğ�PuQ���,]vδI#N�>��y�Y�U�q�iY�
^T~�=Ɣ��j�c�`lB**fU� ��fۜ��h��Si�x|�Dbć�����[CM�+,�g��Z�����M���U]8��2x�NW+�ם�S;���`3~��֨��Y����[7��?_�'�G̞D������gp�?4�J����$Fv�̵�5��������~���+-S�u��%h�J(*��#>iG9&�Q�+v��U_lˉu������z�*�R�h]�:'`���"�%�)[��C��b`�8v}��J\t��*�3z�H�������������_�&z3��B3[���X�,��2Ӗ��9�]�ELQ��)E,�Ie��8�
����7^M9�����/TۆR���$���EYI_M���\L��v������G?
T: ��~�.J�� ��`�K@��A�3օ�iY�샬�:F�C4�(?�`d�_��d���J�k�h�x�D���ya�ٺ馓�_3h�v|U&��A�Z�p�d�n�S��I�-@J��A���<��T��_E�γ�}��1j��b�A�(/��R��o��;�4�i|/H��.\,�v�L=�̵5�\�Y�Һ#X�� ��=/�l���g�Z���k���n�vZbZ���9��d���`���כ�٣��0� k&�୨���ƪ+�6��!��Z�G�Q�`�O��_`���Y$�gŴ0��} �O+
f�I��΀]	�.^e��Z9r�gM�W2Y��@����6�1\�0jO��� ��ԝ��<-ZV�[�I�u����/���Ѿ�Y���!kZ�B�-���d��<�4ү]=� c���p�L��J�����i��..�BՃk��b�A�sf�.\�k	uq����}���2Ķa�u��Ȏ`�v!wA�a7Rc�����/R����g��Q����sS<�D��g{ue��E�z'�l��{t��_ 'E��%`���(ylE5���9DJy1OwQ�>HD��q��[���3̏rD���WK��+��0��nY��AW�j>|�4O=�lRf���e��FTv�^�p�|`�ymK��<�B��U1v�H�X�p�C;߲.�K�Rg%70�oi]�0�ݴ~�Q�`.�M�u=��sD�	��'u�-�tH�Q�ZnG�Z���e�5SHG����<n�И��T��!�$Y�����������~ �ZHC�4A�4s����U��iM�Ձ$�g�o��58��ӓ�^~ǒ@r�q��e��i��G'�991$1���L�Nx��9ԋ:����8���6D�M�"��"Z_�(��6ZqzI��H������Uj�l�i�+h39c��5�c��%�X��.�o������\z���ɴ|�TP��E[���FiPE�E�:�RLt܂�=�������P��yqG���r��qW7���J��ȍ}�] �e>�����FZ��,����2�9��*4������W��q����d#����X~�����hMG�()F+]ֆ��ߒ���I��x�C9l������<�� �Wѩ)�X>��T�j䚸�R�\g]��R�X�Ο�LYz�2�E*y���O��u�|��!��o�m
G��{�cυ,ṥ&A��c��j�������䊠ٕ0ǂ���5\��@�&@b��F��� 4��(�4'�kE/�󵷁��������"[B������[���}�9uZ��
:�)�V��X����fRxٜb�9&Y�G`��U�w�4�5C�c�!7_���xw��9�#����Qŭ��F�Q����7�eJ�8�Wq:�m�2ZӤ5{����t�����"#�8��?cR���T��K��f���0�A�S[��?h���u����[��Hs����x��@�U�8K�PsK�h0�>[�§��,7��\��QQEDK��v����������<̭-��c�l������Gx����V?���������k1	�2nr��6���Ur�^s�\Un��A��ȣ�G.�����-��EW����͒+�1ȯթ�8s� �"�g�_܆�H�Y`�t�sSRJ�?E����Y�`�!��ɘϟD�9+�P�ɱ -�vv�c�ՠpE��3�����?�k�$,��%k]��iDØ".W�:���_{wg���(*��x����m��]��b�����#�v��;�]4D�e����U,j��^O��v��U��p�n�t7�Rw�ƃJ����VBuv��^��I�Ձ��4S�� &�$���i�p�VCy�#�(�5gGY���z�]�����m��ڴ��,������r*�0H�F6D�S�|�8����R�\M���zWP0Qip�??��O:UaZ��P�p@�y����G�R_C�0�@%P�-�U�!�^0�\
0��	�i�}H�*��Γvė=��'0�}Uz�#/oZJT;���I����ܻ�Lv:끷��c�אn@04������!Lq9�߂~X�dM�(X�1�4ץ����0O�3�\&��Ik�z2p��]�m���D4��ޚ1�<=��܁�m�Xl�'�v0%�©	x�}<�5:�tkܸ�N�@��f�������oҞ��y
u��H�J)��Hw����0ץ �xG��2���j���p���(���L�Ex|m��֢V��ݭ��!��ʆy�
W
��Q+�%oa�M8X��V����N�U�bn ��S^Zq����.��vP�'�j�KY�{&n�x]|�ʓ{6lF�s#�n,�/+p�f>,H�)����ci�h?���À�U6�w���_�+ب4qǴ���]0jw �``�M3?b#,�<��� Pq1�Cl<��f��<%'\0�<��uh�)G	�=Ob�/�\v�TH���M�k��y��r����}#�� \�%�˵�����M-�>[XS��fO��l|o8t�E������� }���)
,ӴE����� �Kr��T7��T���
�<���3�H���,ܨ��U#&#Y1;:��ٟ�R�����lxa��$uqǨ�,#v�;_�HC�|�s('7*��_M?�ĖYVh��7�ٛ��E�G^x(&S��.�ߢf�k��P��Lb��˅�M���L�w]SM�U;���O�y�_��Z,�a��w(9����f����h	�[�� <���rl�6���Q�m��Ԩ�h+6'������RyE?�x��D�́�U��)K�hRm�� �+Z���XY�㸥����!�}��A�
��a+b-��\�$�Xd�	N-,s�7�7��T.�L�k��B��b�pA�Ԅ=�g ����Oth�B�V��܁n��m44�����N"�WD��\�L9g���Nk�HEf�G�{�O�u�ZMs(����vl^�`��W��v�}��7]����K����n*�[�h��i���xOL�Fŷ�6��{0Β=���*�v0̇�T����9�Qf��h�u
�Xy�l��N�����E��`������D@�&�p�9��+)�b�X,a�L�yt �����Z�ͻ���˯�r}FAO,.Q�W� �7t�xMGY^��j��{��Sb[�(�_q!N@`O��Q&�W����H]���c�n;�U��.��n�L}$���A�Q���O7�g��:�a�� ����·�74����3�M ���XI�+U��g�R祴XCh9x0� P�<N��g�R�m�W��_lP�Z��꛵ʡ[r�������ICz�[��Q�`�O��]#@hД�N�F��l��L~!��h)��W+��'}��?��qyM<��~t{�nm���S�a�)���r��MN[\��"G���u�v,
�W�/,%�+�P����Ll� ��kBFJT��c��I��W#fQ��8�Z<��7�#=+1K#t��{���7ɡ��.�,�ܲհL��|�f2c���U��r-�u���\ʋ�i0tIln�v.��������ƇJ���P~��q���;�m}�՞P�h�R'��������^sz0��p�{o1��I��1r�@�=���|.����43rN�B�2��Q��8�F�Y�E�vZm��Ι�VzY�	9�!��+�Й���a�i�&�m�ɮ��$�5��F�A�+�"�i���-�<�4ɋ���C��8<� ���>��\�s�˗fu�S�`��d9�*��q㤖�DS[����e5=��B1��``�(t�W��I�����O���������������e.��b��q�+�ޖ�)�%b����|���$4�䔚aW4@��燄�k��9�H9�q�y�-H�5@��U7zN8<�����V�&`��eP���˒W9��]%:n��>�Z�a�G(vVߊc���5Yk�~�-�]{#���o�Dz��"Մk���Y�c���|�K"�[zCfV]FZ")@
O�E�e�o6�B� 6�Z�T�[��~���Sq��7��`�a����v|�}ڨJȏ@ioyO>^ɵ ���rB��W�P�6�oa���~�\��U�����g#>h��ǳXN������nf�(���C)ZFw�,�+��C����D�PƊ�����U蕊�6����\�L�1k%��홼���f#�1 �oe���e�Ĳ3$��iN9������d��u��0G%l��qo�~�vk��ChNXei���L4�(S�ô���j롔3�ZF�+�/ʩ��z+(c��l�[�������ŞW�O�������z�o����G��5VӸM<��O6I>�O$̭��IO@����j^-�
d��Ʃ �Mċ+-�/�(�{
��%G<rOaK�+N��v�1N8"{UvK�J��i�}م� �� �O��w�R���:�h�@�Z�[�|J"�ўM��zG�gWXp�*�D��S�j��\��q�f��9)�lW���~���%�6ڋ�6U��e���z�v/꧲{ N��L�U�a����m�eq�'~�߷m�����U s�����'&��o����ظ��؏Ќ����/��<�\b"D�4G���%��}W�~���<<frtJq;���"P�7bUuz�hAj��r�E9'�4q�t|sg5b���j���l�m�]>�j�"?�f:Zf�CCB増��bN��q�n�P[��_>ӺC�g��Dh��-�=�-��C�S�eyxn��`�ӈ5EZ�p���{+�	<-��ڪr��rZ����N��a�RV[��2k!�=�Z������M�g��+$m�b�F�p�aB��Jb��װ[�)*�`�W����mE��(���	�T�������[��7�U�e �tv?�d��8�Pz%f�^%���X�����|����2��r�9F��R��^��҄^�����B,�bbh΃�5�P���S-[6���|6xi�!}>Pw*ܤ>���9���&�O��z<�ET,�|MB�9��G�fB1������$���,7Ż!���Ɂ���V��&tpjJ6��� ���� taU?����%3����'Z��ƙ�t�x
�L6��Ay�"{�Ǣ�#�?�k���1A8}C���+�lsf#+�?d���xH����燁�ՙ��$c�+�蟎�=��S��I��p>p����]��3��I��!�����,�؁Yh�u�
�Dyp4��>|��B�w��P6�}&d���/���6(� b�\��z���5�X�u�]�%�h�9��.��C�������!޸G�e�m�'��"��+*&����1+'#ò��ۿK��.A�hO:Tae��g�RI)-զ1�%єM<d؜�g>�ll:��o�̅��s-eXej�]�ٓJ�K?�z
<$S�}Քm����#��1����a&���y����է.j���h^cC�֙��?n�ɠ^�Y�#qH���V���q���p�.UOe��,|O�>znpp5��t�Q�e���5$���z2����٪�)�)���ǵ�H��>�\�/��U��p�NxCe����?��ִ��rx���e�]qy4�L��W�nWy|_?�W�����c�2�Y��t�U��m�ƅ���t��`���
��I\݉������-�	������8o��d֖��]N+N���>�{���	�y���\�6~��`����N��^�̮��%�E
B�����IW�Q6.b�&�����~���	s��������A��~��X�9/x��g��U��PEm2yK��&U��G1d��Ę���!�ts=��ܖ3�Ut�cs��X��������q�S�Ib���Jy��I¨]��N�ͱƭ�w&���1�L�k8���K)��_�^����p�3��J�:�(w���xZ �5�#����p�IU���Q�ᒦ{�շΫJ�Bp�TW�>:�Q苖�A�_��@C�b�-Ú���7�Q]�b���\}��ø9p���j����@��R ��2�[��^e� ~$1��R��2?VL�=���A����G��C|�ɘ1���8�PtQ���Ҵ�CƠ֟��m��QH��jY<d�ƴU;��sE/�G� Ɇk��r�� wS���A[�4EiL:s���p�]�Yg�:��Pl S�r����n�O��K0ڸ�H����,���φ���>pԨQ�����7Ab�XfU�D�3�,�����w�l3��%3@���RQ���M$t��j��Kx��^���Ǧʠ"�魐O�ߙ�!�X���l�ڙMJqG��+�,�!їӏ���2V"4���:B��ZŹ�.?W���T��ʫ� �Pkۨ+�k�Y�a��IЕ,��X9�m�KSv5qӧ��`Dh,��g��7˶)�R�֩vSi����]Sa������Ds�3Jp}��������k�"G�P��Ƭ~�T^iǦأtҰԠr��`46#�.M�ܶ��Sۋ^�^ĵ?;|�u��Q�P�cyz����L[��b�y�C�D�4b�W�O�lQ���O�d�h�o8���ӻ���<������AN5���p����n�#c�|�+���:��N� r�o�`�
tB$�23ycN)��5�@��v[b�p)�V����3s�`�����a>M׈tE�Hu|'�����J�qE6��d(�ʩ��-�ڦ6|���[��W�'~$�-�a����&AIQ>�������Z��x��Vy�G��oK��C�WpZ�P��4�Ug�-�+�Y4Q�SG��Ð(�u�)��ӡW^��˦@u.����O�a�����9yjn'!�#O���T#� `�u��mq��a��fo@E�O����������5ěy��k,�?Y]T'+@��E�%9���p�/œ3�w1�����rc����G��}�D�HPD�KN��i���`	�nE-舌�;�� �'"��/~n�l�o�ךsŨs��%9����b�w-$�]��
1>k�I��l��$����߆-
geNШ�e@��O�_}�[�\�P))},c��s�TvPOv��rՃsh��5��n�a�Ƌ�+g��X��~Z�kus������	����am��g���hb�.��i�ˏ0�9���"�Rvm�����c����R���ڇ��"Ϻf��t	ڙRf�q
&JQ2:(,r��4�e��'b�s���Pl��S���t	���6e��Ȕ7m"���^�S^��w_�_/��~����Պ�+�f=�७�u4+�
XU$o�ӳ�y}˩������}��A��C_�9�h��`�o�PA[3RU��I����Ⱥ��ѥ���]%p�������}���Zn�;�P$*�DtQ�9�[��"��<�/~Cf3�n��,L	�Õd� E�1��g&#�}�((���ʋ-��2΂Vi�t<3(�[PY6��>(v��h%�$�Ǿ�V׆�~�3��0�m �y�`\� ��E'6�]e���aa�R�n�N�>S=�+� wyD�L��AM;�����>^������%�O��<���fy�g3"m\��Fʑd�0i��Y�E&_��A-�������H�c��$Q2S��0�-�ũ��z�ͦMdO���6y�A��	�i�����i��>4�L��Խ"�Z0k�q=�%�Wo4���ɕ'����%�����w�G�����������F7?_C�hЫ�QE=sĆ��H��RT�QK�z8>��|'݌`�S�	�Wj�D�+NN��O����bG6���(y��F��߸[j��
��҅���5���P.f��5p�E��F*��?�����K4O�B�������i���\�'/x�#�n�B<]�7B���^r�be�g����;��i��E�&Kګ
�'%�^9���_h$+#aLB�O�0�@& �&)_����5���Q)�8�|�S�4v�}]�I�E��M[����*����E��]�t��dkb�`eC\	]
l�i�;�����*@���HZ��R;FQT�7�C�~�`MȠ:��:noٖ]�/��QY陹
�QJ�(����"�/� ��s��J�`r����0vf�ܫ��P���ǯ@]�wj�CAO^`�Om۬�z��?'T&�)B��	\=�h2}�N�ϣ��z̾�L�����B�|�/-�M���a����vm!����@����́\�S�Ҏ�� ,α�:hlb�ٗ�ٽ��e� 7H��T�y���NAP�j؟p��"�o5���\�5�\�e��Z�4�N1d�!ՠ0�������s@��.�0i�j���!e����5�gA����G9�`W�	 �sd< �f%�Z����G=��]R�b,0�Jk��O����=����?<�{�-Ԍ�Sڐ�F��:Y������x�k!oX���n9mp�f����{$>C@n�P�P�ɭD1z\@&��Z���OuZ(Y̱�^���{�KsWe���3,�~�rj~љJ�,��f��h�|�ќ�%ڃ�@�h'O�a�6��ɕht�L�I��g�ؔ/���о�B�ǣ/��$�pb�D��B3�7G<a�4��'y��#���=��: ��L�g�!,-W�����N�M��n�D�����p�V�]��&��1{�4;h�tV	�e@����[�D-�WEn�W�K���;�������J�^�Nn9��}q���e�����9W�u�#��n�o'gܮC?�W������l��//�J�c�9�uNF��;VvG�!��7+*�!��R'��<�kWH��3�ҏ%m��F�z+~6��݆����>�4�A�T�y��v�y��:Yx2����6щD�&�@5�x�I�,ʄ �\;��c�0�h�^,(�Fth����%�`��V�9�=iS͹N�E�|��p/�yq0�����)/�����O�ؓ�\�a+D�;���Re<����v? \��a؛�v_��J�h�O��@�I���!��i�R�Hp��W¤�2��{�� �d�qJ�i�z�%��bfq��K�q@�с�Nz7�ً��ˬ����e9��xūG%�@��ܲ�j� 5��CG���@�j#ʃ�
Qb���?%ޱ>y}ȫA�u�7�H�nt=v����!���P/�:�q��'�Z+�[;��x-�Obh5��o�?���U����XB�,�D����cȊ6�`�����̈́�u1^�9�<Mn�Bs�{�m>��އl�y�Ɩ(sTv-�~�]��,6g��»���s%\Z�k�4wԏ4�e�7-w�+;k������b� ���p?����(y��D�]׳Y��\��y�S�;�a�Ui�]l����h�L�H�	')�0�\��VT��Η!w�共����<-M�Ն�D�R�t�.>��k �����V5c�a��m�<��N��c4&J{}��CP8�H|�X�	ЎQK����ip�dVS�{��8G�L�?�׽�~-��!ǿ�	\����H�h�t8�����}��)�)�����o͂�Y"���EKN�m���龽�V�3/˪��3q���x�j.�\a�|'6 �Fz�Jf���� i�\��W!c�?��g���2��^�q�z���(�t|���d'}�n09;cy7Eʎ�棖�K�s����b�^Iv���3j�Ҽ.�5|�2���xt���f�AY(�`���Xs*�����߸@_u��R�y���[��\�Ӗ�b2ctSߜ�I</{J�9�L"q��J`Sy���4��v�Ņ����\| m��;�R'8O2�:pP.��[R�o�R�t��K�Y!��\�ݼ=�>�8���a��)f4�n������{P�Q�Z
��>�2XGD��p�fv?*� (,�"��i�����yI�?l��0  ݑ<�$;��>�p��\	v5O�8�0p\WH�'/d	*2������ٯ�Q���b�p���Ϣ�������|A�I_ŗ{j���ܳl��k�,���� �N^�+���w������{h��~�q�'�A2um����;�֊'�v�k"�Zg������'��H,ɑC�{�nf`���6es!������j�����Ig�ʺ���SϾ�4h�l;[g`A�z��N�lR���s�~�䇪S篇���RK>�D��z�Ƣ� sr>>��g�iΖ��ޡ��������c$�d���/�qo4����7�7,���d���YV�ށ��RR��XܳN/J�4���9Ԟz?��K�Ȩ��(}�K��4���s�y���	�d���I�R�U]SdWx ��l����I�'�K$��iʪ�fؠ�s�p�yAG��J\|����Mc�n#M�� ��qYO�p��6�)�[1��~�	VߠP7r�(�?J;��������Ҭ/�����W�'	�/���I��������F�_���I>�����O1|�Q���	��8HCK��p����)Q��˒ക�4ళW�<��!?�����	���Sitb`K5ߴMm��t(/���VjQe=�����/�w(�������3���9�G�s�A(�G��~�������^2��o_��8��D:�b{���]���2l���[���K��=f�w�TJ�c^ �ᨫ^ed�rm����ḟ�OR���%Z��QG�E���><>%�-��c�s���S�|Ƌw��.����m��R��n�u�|����H��'����r<H���p���T:��E��k���� �~Z�w1<D���`�	�[n�t[����-;��xC"0w?�������ll��(D���ń�I^a9�J��&���Hj�� ��%��j��Nq�#����/.��Vj�K�`?H�F��9�d]�4\%��Q������p�K�=)D�gUd�&���+���Ԟ�ص���L	��a������y��ʕ�)
`��P�4��@W�0���P,|�ʛ�-%k�W+�7ǰ#�K�h!�1��g�%0�\�P. cn'��w5����C1+�v�>����p�|]�~����V�D�����^T꾷��)/��<�c=�� ��0�L�� *t@�OǬ�*�F��<�a���������������̑��J@ �D _Z$��77?>��t��֮�%'��~b������o_��bOӨ �5j�J��ԈT�J1�'��fw�uUz�03)Bo$f9�3r��1z�	H4OW�T!�jc\�F��'��<��w�������3���)�v�ebn��sNh �AP���&�دXfT)�������,u<!4LG �����Q��ݰ�qO�TNG �y���bU&׸\�ȟ�3U��PC�� d�^�]����ZJ�����&z���*u:��q_|�i��Pё#d���z��X��V����~��Fe$�9��?����"�"d��w���W�kz
��k%,��A92��^���ֵ�?���]m�IOy��8���G��|����;�����y@;$p��T���d��m�6 Pӵ��J翘`;]��
�td��W�-��y��K�o@�r�pYkE�C�dBqq���_�zp
�b}�l��j%�(���������w:c=Y�γ��W���
���{�5
w�kW��d)N��]�j���Rd�~��0b
�/�Xw[@TRon�˷|��^$x�J���'�jxc���y�g=���HD���ƒ
c�*��$�F�D���C��I��ġ�$�	�j�K�(NW+8=��FkO�cbï��:��)+�53�Lj��Yh�.J�A�B��@��0=e����q�����^���$�hQ�a�-ixp��QS,�q��4�?Z���� �Ƴ d.:d:|�4T��Et�f�q�4�"P@��|]��w�/��3�E�ǋ��]�H�j�8�M_�:x|��.�b���hCF�����&?`�4�Ьe��_͘�`o�^Y�N5�"j��@�h���!�JD\����2b[9.}��6h��=�p��@�y�FP��s��D�>�AxdBn�;��*��m�B�T:'ŷ$8M9p������K ��ܔf%�n��L���{�&�7k�/`��֧a]�򞏱�^�����Z�U����\��l�Dr
���#����,tl	�2���5�Xk�3w���^:�K��������!�Z���R��n�*�G�(A�8���+�e�G��"W��HI��p�_�H8N��C�<Jsv�ݍ�__:��¹����aO��>�I�8Q�9�S�7ܡ���vl���M�^�G���`��An%�&J���U��w�:�xʜAgg.'��2�N�vEd��� KǾ~)Q��Zęߗ���7��m?*�8`ӷzJc/ �uG�i`��_t&RB1�ɠ:���dB��	u+���fJ�F��F�Ǆ��ק}0��4��d��x�S��}D����ܕ�~�.��V�[����)2�P�c�O����-��u��R�]�z�kD�s��A��ۤn��ܼ;Z~G�=���d�zꕷ�~������	RmXCi.�a�O��!�U��fk�i���xv�����?�������3���A���ѧm���բ73OM�:��n Rsr�����Zq��!q��j!!�TB�j����!�J1����zewA�
*"}��jp囙?h��[-쯼�g�p�G�K2gq_ֵi�.�a�C���[1!���V`W(M�v��EC�Z(F3�QNt�$'�_�oۤ!d��\�Ҡ���D��ox����[ZP���&j��_ �V¢y�x�3]����"o� g����אcX�Xz� ���K�b��ZsT�b��㇕��L�lA�#"y���r��g��.L�~�B�j�L�L7�C(Y�y�zcibA�}��4j�G��1�(x��������)~�n�&h�=Jx�ˤ�ܑ1�R�����#4<**��&l(��N��ؿ��[��v��i2!�u�ɪb����c�2m��r��kͤT���e1S�9xw02��YQw�:�D�=��Cȿu��oU���Q۞�S�59�s�3�n�ok��Is��c���7O��k�,d�>S����-��;1.�z����佒�{���,�Z�-��u#ZJz��1�g�58y�!��R�I^�R	p(�k}3�t�I��:�[�^j �aծ�D�*�|���\�_�XV雲��`����a���KcǰY�lU����aB �b~��Gh0|�h��(I04��2�;�حa=��ƇC[��}���3o�Cz�Y����-D+y2�P��N������/ I20#�$�_Ǒ�����4��_��z��Ĭލm��dزS�b0Bc�hñ��Tr�oK�3^	�e���J��R0`�澶'�4��{�����g9�N
�Ƭ��0BҘc��օ5��>ߗ��=����?����&@�[l	겟�DM@�� I����1�K۝�Ѯ�}{�j~xb��x�>�y���+|�l�7~�����0�IvH1r�1����3p}M~jd��ڵG3.���0���{��r5��N0C�+��;Y��̪/���Z�Vf"3b�fQ<#[d颎z���+v��rx
�װ(��6::��j�:?��H���gT�h�B��j�(/�%��t��]ж:�i����N��Mx��'���6�}���U���_cA�Lk}Կ}�+��N�J�g�	1�G�nZ��N��H��[3�I�e֥oa�������T�ǐ|<�����6R9��ϰVD��0|\�\�j}op���YBh�QC�U�j4_. x-X):���Qjow�^�p��iE����^z>��[�a�h�!ɼ~��J��M��V)/ц�ւ��h��HE�j4�
�
���f�+7������g�A���t��M�Rii��a��uJ0�k�����ʈ��W|�Ə���o�,� %�����{���'.�S���Ҝ���}���I�yg7��E~�}8�^`re1��z=t�ӏ�G�˸��J�C�ݫ�ƌ��ϩ7�;ӺR��:�cU����x��p�P@Z)Ɣ_8~��?�N�0s�H�g�6�r�Vd�p��-@��ʥ	b.-��Q=�3q�S�!����!�T�SV�_�u�%����p jAU�#i"�X������b��gv��_�Y�nԪRd��������0��5�ԡj���Te�
Y�(D� �����#_N� U|b�%F^�or,am9V$lr�7+e�I�h�P_\��gQ��h�eUWc�ǺU?��St(�_ށ*J��U��Ed?b��\m�M�n��#% 	Llw3��Дz���7q]@y�%�o��A��&>�VZ!��!E��V��(�}�9Y�r�{f�� �ҕ���ve��}`:z4���r�lnh�R�,b�	kY'f�ί��b�U�xz͗c���ȌR����ô�i�u����7��9�ûU�?�w]�eP���g�I�o�v(w@�E4cs���]a��|��R}/6n��5�2t׬I���D����[��K�C�X��N�*�&����Q���W�}��MեT���wղ٨e3-ˣ�����4��� �����:	'�*��#�NO�1����˱��T�SI���w��|�MI37���Ԓ�h��_D��q�F����I��_ۏ­�Xl�`?A�T�I���ߌ�W��k��%ƩK?*|ǳM��M����j�����u�~���� �;"T�U���,n�R!ѧ���5�S6�$9|L���/</֎���H��k����H��^r8fD!���0R
:��)�8v���?M0D0�u�IR�7~���pe��Y��L��hXD�ú�uŁBC~�����D���O���%0��Q(�������n]k�h�{Q���;.6̽Kp~��	�q�[�M� ̳ �+yݯ����>`����-�k��Zq#\^��Ɉn�o/��}���-��M��6p��;��L�q�Y����&�wM;)p�*$ D��hW�?iέ%ۣ�>��A%��U֋Aȓ�����f+�',,��7�t�!ܣsi��T[�W@�/����M��f���\f�@�ZL�!X���K6���o���`�U�o�1������7���<~�k�SSP�`6WF������]���ᰃ�&��L�]�f��	����㨗�I�
׮�����YW~�<#z�~M\"f?r���,���i�*�Rl4��FdN�����H)s��&�ړ} �0�O��cO&��]z�\0����%l3I�X�bh�����!.��\��Z�zr��a�F�Lo�t���k3u{Z�Ђ3m���=@�1ah��^XϊA�D�
�L��(��	�-3�T�C�`�w ���^�)$�>Y�'���^��K�SjB�
d3ڌ��6M����L����9�v �/қ5OJ�.[�B�A�Y�T�-sAqV����y��/�Dl��yLJ����ele�A�D.�Y�����%�A���[���'��zk��׌�D�V�Q�<��`�,��Q����PnW���U[�8��I
p�)r�(Y`Y9�����*}׷Wj#n9:��n��(Ga l�x'�)Ä�6��� ���H[��N�Į!��=Sa?�/.i���&C���;���a��Bڦ��ܮ�bj�����������:7�#X�ːyǜ�i졃�]^��!�0�Yu�I�NBs���#�ϫ�H�E΅¨��
{~���6�eb�N?��&�Z5=�ŏ����2�fD��@e՞�m#�)�G=��7܈J9{�<�(���G~��Zd�.�M�Qk	*3�SK�ޢ�� �W�B��jW���N�W�8�]F�:'j���wf �h�C��ג���h	Y5T3����p��pQՂ.��ܬ���8u
�l�<�����,K^�L>&������k?��1)s�6��>�4�^z���k,+;�k�?d��0F0����H��K�Ѕd���E*T�'8����v�(�m��P��,c�DR%��8Nt${���Ye�)����q�G��:��"&��&|�9	2��^
/���l�x����~Q��o+u�E�	�4�\��Т���j��[���o�*+]t���o�:�n�~2�ҲXz�ʱ-��8_H����銦i�4d��;��:�&�rzJɔ��nne�:�;�.�=h��!#1���$��i�T�_�A�����k� JU(fO�-P�~����Pc��#�fG@fd�ut�V��"��N����Ab|�`�͙#�D[��R\�4� ��}��8YA.���O|'r��ç�*�*)�IS�k�*V=�E 3�p������H��>ahU��Z�q2�yv�#դ���C�Ъe���X��5{�В�wė�E���1���ݼ�Pc��qY%���Ǝo?Aza�͝y��d/'�[W�����]��>���瘦��h���hG�Nr�(� ��%Wz����_4��Bu{c0��漂oP���gBrYq���Y�F�'B]nO�$l(���c����"�e|���\f���E���dN���Z�����^�� �--1�>L��s����]���L����`z} P$��`��R����4-U��e�C�[�fau�Ϗ�������|pR�1ɻ)D#cN]]�Q��[��0ܪ���5֐v,ը2�=���ln�������m�cUm��{�+op�h4���&����FL��E��p.'��5V��aR��� �9���w���U2�xq?[!!�����@��٪�-9���#I�¦_HDM
�-����ټ%����/��=����5�p�
d�0Ԟ�~+�f�~v3�,�p��Q��
�`���O��jď�ْO�0$�D]/����	68�,h��|ݥG�o�7�Q�U�ׅ]��.�Xw�2���{G�� �vWu:)d���|��x
}�";/;��u�|d��>����߲V�]̮w�Y�OV�kj!O�[�@|�����	>�<Ȃ���n�L�RE[랞�^�3O5�?Y}����#�{��s-��/�}2N���~G��0\7� \��g�7��Ί��B�'�N"gf�d��Cܞ�_a��c�:Q�툘�T����l[�bn�lXnU|UW�(=M�W�6R��|��5B�"�﫣�-m[��u|޷�oH'=�Ɨ�-��1���Ix�g����`7_e� �'��ܞخ���-jnJky���œU2���/�}n�27����n���#6�c�$%ۼ���^8QW@�XG���N��G����F�U@]@���1F�(`X����jn3���E-���[��M�ʗ����=>�S]A9W�j�T*=��vx��HlOȌ�o��a�)Q+J/"�U2�=�=�O�b���C����=��3��"��0�r�>2���k��(<� �
[;�72�yУ5x�G�4+A&zY�l�/� ����wa���6��UN�`}�J����Z���y�1�~���ҤV�� |�
k.�<U�yĆ�p��=����!��ط��,P2�f���*6����#��ү���l,v�`j���3 O  ��#�*y���=;Wm������ܵX��t�7Q�r�y�N�\�=�j�^����R���L��1L�i_��q��(�H�kf�
�N�q�ی�[^e9��{��Ϊ�P�e-dңݛxpN���Q��S ��O�ƢYy�)|XǒQ��癬{�>5g��x��j�}�X����m/�S�[k�����je8�,���[����1y����o�N|X2%�֗��Ĭ&���"G<V�/i��?-$��;�y���<�W#�O}1�
�Y+;"�ٛ�pMRLbS�N�덃��S4��@P�Iuj`׋x준c,
ɯ���n^��1n���4*�G�w�f{NZH�_����fi1Lզ6��u1‥��{z����Z�7���NQ@R�� 31'\k<׵s�a�4�n' ��I�V��AD�2��Io;�����(���]UV:=mU<��S";)̄����pR��+� �LNKv;c~+��1�ڋ�-#x�8�
M���*��]�@���"q(kB�V�r�6���/�JM���)s�P�l1�,�q�&�p��A4	't2�\"z��U+m�9�CC�;�_�z��-T3Ϝ�ԛh�.��,Z����7K���j?��zL����n��d�h{��}��D	Hα�,+��e�.���|�����nހK�/��{��`?��E>u|q�(���7�W�.����FC��'����sH�<�O�����d��G���ʧ���~!\x�h[G�3>U�v�1&iT�R�C�����E�K������#�t�!+W!�Pe"E >У m���ZF+a�G�/�,�	k��j �����z�-���W{�'���<Ӎ��r�H��i3��ͧ����2
o}}k��vTNm)s����[��;����Ȣ��U/ki�!� +��� "J�ƫ=���젾 z�D�����:bZ���l^���0�ԃ'a�֔��nu>���b�M3i�,�J{S	�f����!D59D3�?S�M�����{����w��l�iҩG�����3q��zg'��=���������U%?Ͱ���f&�(�=�K�[L!���j��e��r�����7��z��D��F%-����3��*�/|R��<Y��	���Mn�����b�?�n�]�+�9��k8�1{�d�
]������]��'�리�g�e)��f�(���F�M{|�k����Kb*̬�������<�bN���S�:e���4\�nC)&�������<ҿ գ�`nM�]��M^S-DS,��oF��厌@7��ր��P]��Br�>��mYd� ,���ò~�{���vΫ��G�H�AvlZ��$3_s`�~$�:����@�n�{q��Pn�:���֛��Z���d8t�7����Nܰ2��	�	�e�&�鯀���-�}�äw�F@i�iC�_���v����k�ޠ��s$K{���nqPG�%�(�,�(.'���!fo&�+{�\�Y���Æy�[h���Jo���$>l+E�F���!')5�C�G��]hg����=�燐���cx��>�����)_[ G��.6�l/�F��[[b���|�`qH��Q�B�}��%K�`��3ާO�P	�"|H6�����]��H��=�LD��*k�6��B4�@Jt��|�{u���c�b{�?���e�?���4��[��
��/6��dc�݉�Q6�ml��Ϫl�=�h��>�Yx����* S1��6YL�����6��YگO������0��b�ϭzG61w\^^����u�'Jކ��.���i� ɡ�4r�
���b`�2.��ʅwJ-�V�W��@�������Q;e��򠡪{uHo�^�AȐ���S�䴶q���=8�ZM
%9 /�pԢ�) c:��qD�C6���"��X���i^�����Qfv�i݂w�P��{���9+�fۓv�Qd)�
�ڈ"T� �(o��bx��s��&��cN�|I�ީ��w��p�TA�:��-֖#������|�-)Z����%���Q�[ɝ�8�eB���V�MM#(� ���S䚛&sk\Ž[4\�K�.��f�w����=�>R`��T��y���n���]�dN��� Q3XEp7nn�jӠ�ll�O�T�W��g�$PSU�g��
�Pb�`���^8�k���=ch�,͓�i���m�� ꗛ� ���X�"53�N�.$�E�Mw�2C=��T*�'G�oU��II�	�J�K��3[f8�u~gZ:���H(��ا5�iu�;��ȷ���p)j�G]W�?��`Xr �+_v���*�M#&-H4h�����(	�L?��(��(w��H䧱���qE�i�Yfm>�.�_���ܐQ��T=�(��Z��I�۴s��/�3r{�"@wڦ�P89����P�M��ƶ�9�I���ƤH��G9�?���͇؆1.#�"1�qހ���O���CE[Nq(�����n�M��>� �8w����MP�?ᰚ����$��Ǵ`;���������L������QN��"�e���Ә��|wx9|����6�-s�	�~�ڦ$@Z�|dP8Z�B���d�'�)Hu�Vt�y�Q�஠Q�Zp&v����h��r1��4��oq�ا��pۀto<��z��S��4"�/-ow`![�hWCS�|�����vV�&7�7t*�l$_�.�����F����Q�x�/���R��J�Ou����xh�^��4>���
�F�@�4��^��F���jL�=�Ԋ6���ۑ�k�u�4����pm��m��'Ǒ�d"V�ł2�p����|�Jvh!|ٙ_��!��r��X�6������[{��:����&[�!�Yfv�M씱�s�j�wY&��m �A��Z�e���Hh6���^l�_G�!w���n	9�C���k5�~ͻ��{�p�,�A�N!�dˆ�hâ��7wvrok��
�b����dW/�����Q�y�	� 	oo#'ˆ��6���I%����pHU�Tύix98���ja(,����#���ug��W�o0��"3(2	���	����V$0�ZB��������e�;��[��z��ݨChCg�f�Ms�Z��Y�̞�����F^��qF�+G�\�*��C�=���{��Y������t�Q�c��v��d �7���N���֎x6}��ﬆ�h��a[�NW*��*���U@��~��U#d��j
�؆a��&��5 qy	��h�BK�4_�R�*��M�Q:"������Z����\y�\�Vc�-��;�������w�w&�kϫR�����%��r'�S!�1����k{5�:#��W�C�x��OWX�H����,�xq���t�
�ެ�Ë�������AG]q$��N<R�3�ќ'�{�v�T�`ޮ��A��^G�Q2<;*x�|^6���� uk���fHP�W������:`���y���成�Q�z԰�Ֆ����ERh育�-Y��mC�F�f'���̐ʸc,��B���?�f;���kV_�����&��o���_}WC�Q��L�Gt����H��-˼�QA�۳R���y:��,F�+s�z�
_��楴_F��@.ˆ�R|<�=t$'�����N/��J��b *�a�?�%t�	�o-JH����^<~
k��M����ˁY��p�v&RQq�� BnK����l�O-�Y��]A�t��cﻌ����D�տz�d��ɂq�N��B	E���g&O��?`@�o7/�u��(+=�AY^� ���q"���ù6���I˯pW�1(���5ݥD2WxR߇l���N�gcx�:�n�m,#����Y���h*>fۚ~�J�2d��N�����fx��<?�x<FL���M�{qc{ߞB�x�E�-���?��nD�k�٠�\�����N��2˘�?��c�*#GEC�;�,�^yh�A����\�5I�7�U��� �hw�{,�`���i�6x
�)&|ٵ����6���x���e���@V�6�����ld�V���3ސ��t�S0�ӉSx�D��~t������StHy�E�x!�}���;�1~�h��rw���tj���̔����j�؄<���OfG���<��8�,����Ҷק�1����9OX�1'�K,���l;�\ڞ.�X/��zo�e%��z��yi��5{Q��8l.���k�-�~��f�J�-P���e�&:�F�� �����v/=?�*��t,�̔�Ԧ��2�xNm��^�*#B�֨A�IS=�ۙ��宫��lӲ]��nÈ�"Պ[�Ab���.�1Ќ��dg�[�{K�:I�tk��	��ߣi��n��ڡ���Hu��C9��*���\��ֆ����tZ܇k!#�xWPm�Y{�tL�3�%�(vg ��J�d��uO�K ⚻��0J�I��)���������>\O��.�Gpu��O$N����X̮��"��GSAB�;���GI�C���?����>"�`#'G�Ug���8vѨT�B���V�7\0 �B����?�5�1�I�y�Ԩ��
~]�'��M�j!㫅�7��p	��uG�X`�;ufQ����żO(��P����A�϶F[�I1&��G�a�p� NWx&6_|d7��Z쫎N�h�}Gd�XSzm�!��$C�t�~��K=���{fI3��j��]�l��oZ"[fw ���:ߍ��(U��z�N+����������_��!�D�t2?�Ĝk�r�;<��a-f	#��R`�6�y�[\W� �Ф5�ХقQt�H2c6�Q-�vs�ՒB�'��ӹA,��P���t��2���j��wY���.~�V���t��{C՜�\��!���g��;��T�hlIS݌�LMz�y.cn��?�>��(k��\(�?l�]8����Ш��^&��%�p��.�����E�5d�����j��?&�tE�s�Őt X�0�������r�Œ|�aI2�v,���|�w�D��z?I}�@��ݶ�8�8ȿ	Bѳa�%1Lbk���{����?H�B�oۥ�zJ4FT@��Ocm��sU�ث/B.�5�$q6�{�{I��T'ܨ�?�$nK.�I��#�r����w_���.Q$��3��$N��ڛa�fK۬:�z3:�#�s�}}q#�M�����*/�G��{Q��Hg��Qf�v��"�*#��+xX�`{U���B��(�hq�ȷ������-<��W�GPf[�L%@kާ�7��u�(�C��j��4�G��iF-&��+�tV��[iV������#ga�
����K97������Kr�L,�xBA���:�_��֠UG����1�FG웡hXx���kʆ�M˪�&S08~��Kf�s7�"��-��4<}EȢ���L���� k̬z�CT�/�Ѝ(=�W?P�4�ʕ�bXۢ_�(����zB`�����w �a�em�DQ垰?�Ő���wGM��v0c��;�@��C��G	��!L�]��k��w��K�_zBɘ��_\�1���G~�X+%V��ʟ������V�V�C�X�d�/{�F�r4�~8H.ÎX湯AKX�k�Mc���!�ں���F���e��V��;�N��Pc��g,�$��+��F�}���9�:���p�~�+������?�z�͵a̠�
� �9O��v,�>�S����� ͧ>�8#@\���R����徨;�Ψ5ޮh�k�}�kޠ����ər�7�yW���!�٠�d������T��%�h(�?>�A,��gU+������~�=c{���ԷJ�E$��FRB���ܧu�I�{�C��-�G����si�2�X<��PD�;8�Iֱ�ly�p����ڹ�Hʞ��@ֆ�Wh��u&j/v"��|^si$��-�܀�Bv�~j������~�v���c������v�mMx����|�d���~G�6`�CdC^6�����~>�����l9����_�P^l�g�'.O`��e�2�qH��IF�.7֟��
��i�GT�_��[��u���tCA7�kH��;��:���/`�QL�� ��y С��ro�Z�I�A����)Z
�6|)lShG�VxK�)�Of�:v��C;ߑ=��J�I�����!CԻ^�]�}��4d?�+8�Zߘ��uk�Bw
r����U���1M�v�F�;07�)}���>��PE*�
$�y��`������rCdsW".}ffYZ���pQ�KX&�"��`c�Pg?�f�����=y��	:}�������D��pct��F��6f�8W����a>�kp������KL��ɓ�ݳ�^:m_��C>�� }P�.�tt-�P7�bʞ.���b����߫�J���l������kî�$n4Z� A�n�����m4Q��]�0Q.�V�Pb菹>��:�tMj}YN�'����־X�;�=��uP�ڲ�	ܹa�c�H�;;P��][v�}���	i��n?��i��Kj$R��ȽL��䢳��Gf�ٚd�F�ާ�Aڗ�tM�*<�{��s�w�J"w�M�%�޻�A^Ik�'�rL`��*��Y�lҒ
IA�|�WFqw���~�p��(�9�Ţ�p�t�o�z�2C�5Gs��m㴿�g�v\K�n <>���7i�����knQ��s:�߇����%۪@9jC�CTQ���H�[�&�#6N���������=\��B�'��p��b�!���(��u�O���/��V�V$�m-�p�l[wa���c�@�0P���Ni�쏶1U3w���MW�B��tr�L���vXGY���[�_�`,)mdFRz��;}[Æ<��K��LΒ ��	���j:�����P���2��A#}X��MO�tD�D	�F%�{+HsG���Ue�z
�����[�`x��ph�\.Y�4v��g:ܿ���W�g4?d�;Ho�E�[��π�X���$w��qH���k�~x����B�
��*k/��U�%��%�פ���&x)�`����'��*x4mq�1�<\� :���T�=�'Lu���pGLq�j�W@/-�'��z+�������C%���l�yFi�I1��Z$�`<�>p��G�f6lETm}m-Ms{a���~Cj!a\J�6��l=�	Q'��"DB���-u�����}��t�m�)�_�Q��8�2�[�#� e{>�H�g�2m?L=�BɄ�@�a����b9�]�	��
7I�쉓Dw�dߎ�,*)H�X��.�+V����ԠU�� c���P�=��Y��*ɰ�~7H���ˎH�����{n&Y������~����]�<�y�@����Ǚ�
-�A2L���vW"�X#5
r���)a��l��GXj�G�Dr�a�`4Gѹc��џO-K���%�Z_��_Pۀ����.=�(^};q��y��Eg�񲓡���(�t�2��o3�ځօ� &yᷗ�)=m���A�&*Q��1�[[�M�#!Ԏ��.�w��� �΄�ď~�:RXA<r�?vڮ^4�<���4�Br������TwP_?$Q'�tS��B��򄰛���0�9��S0�)�Vȏ�޺�#�PԸNZp�Q�W����)*�ƪͩ$�x��m]>�Ӱ4�)�{?��zP���F����(kh�A�֡��ԗy�w�Y�$HW�:-�}Mn�y�\l;���Zl^u���Ή�O�Dk.מ��yu�6E��Nݐ����2����=c����{�=TYef<YV�)�?9im����2|�z'�Jce���bV�!^I��>��)�,EF�[9J���+���	;���A��Цuu��
���U#���2�)!x�!ڷ�N��zlr:�*AI:��Z����s���i���0��u��ߛTP^�ȻF�*R��s�!��E@C)=�!r�S�V���L��c (����;�;S@gFSԃ�Q�rŽ@f�[���-���f�����S�����CMV�"tI����،���}�G�K-���9���_4�B�Z�p׍B�B:;��p,�_:/���L��c>G\~������&���!8m��yM����B����	4�l�������\�ĥ
l,��ȣ�3��*MY�Ԩxg3��,�7;����M��L��GN�';//�r�"�WE��A.� R����j��l#��z���4ў��鯠�@\b��V�h�+��c�� ��}Ἀ��5�����>GNℯ&����S֠ݑ,d��dhO���G����G������˂˒"U|�ʠ��x(P�{I:z�.��{�G֒�tEBލ�.�!��/��٘hof:\P9��H��̘n��C��	�5��F:d�ET��7N��El�ɨE��8}P��<�� �w��"�R�lN���O�##�Mb%�q(���ኃ@ov��6��bm�!�-n�
%R;ʸ4���(T+�4�?EB@�j��WDs}��P���إ�Ʀ=jž�վ([,y�Hv{��~���{���ۑ�3��)������
�
����+�jJ\λ���D�L�"��flp�G��
���,v�c6{޴]м�)��#�(�z��ݬ�̪З��DK|�X���]�۪�lrS�L��SN2	Ԝ	`�>c����8��'·�9��"
���mX��a`�A�Ԫ�@F��`-F.2+������I�������ݭ?��mX/0s�7�%B�Ҷ*�S�" J&!^��8X�]�U��vO����at�m;�Eo"8��a��L�0�в�N{��)����>>�F�-f���V�91eۑ�=��&����XҤ�iN(�����G�&�� PŦ<��iB��(v�����T�|�	>v�z�Ǉ5K�
gW�G�g��p���u�`#�]!�+>?oN�c�ǃ~tL%S�Q&�/�5`%���Y&p����7���EH��O�Q��=���f�>�Q�9�Ν{@�'���r������}6S?x���`��LXC���ۑw��'}����t�}�z�'���R�r�Y,o9"4��1���}��sV�&���1����aC�Q��J�=��i!P^uH�e�W�p���WF�zO�����B�*RcE�����U<~����)�Q�Gm��U��@Xea����=땙��MrB�rSȞR���Q��A%��FR>h�~jǼ]wj���~�V�)�
(�g���Y�K�V
�X��$Ak���)�Q\Jg���pE�3._�F�ļ��raS�|���QLR�N��km[}V(�{%����L�l���1��f��-��͊#��J���O�S�
��,�}2�%M�̙���]��q��i�{A$Qk�'�x������I���Ab�	�L��G��G��#?�:�ܻ@���Ģ�2�fݗ��7����82�Lʪ��ų��7�	K<�
M��s
v�p3��7�_n27~L�s���yT�r|�Y(Cp�^_�X�M��	��˫��m�����3hb����q��(��MA�0�Z�C��1;�����\o�ւ~��ƹ@;s��F�V��Sﲕ�J�F�bp-	<�x�q.����\'B����C$�1(S|o�y��aɬC�eK��T�΀��:,�c�rM�ղ�u�l�<�&wQЎ�*��G�["2���-�܏�go�UC(���1Z�Q�*�H����l�^�W�$o��D`L"�����0ϓg���Y7r���o}�|��!%����k0�䙊�<�֘
��΁[e٧T%���_��E�ʎ�Q"���n�$�� ��I�o�T�H����*Y�%+��UB#�K�ٕ��5,�/n`R�����QD0�����k�\���H�w&���{ge�O6�H�Z�� �sR6��a�Y�;���ھ��n(p��������t�8>@O���]��|��0y�C=�;0�)�V��O�E���?� ��	�X��:�3�(��sm���f
3g�F�
�^�����VRq���qϹT�0R�)�P����(9"��Qm�P	��jT>�s�i��3W~SX�$�ٹ���oc���3
����@��dNJ��(.?#��s���,K���o��aS͖+�6|Fj�!akH���C��8B>V.�|�1gn��	֜��a�:�YLhU���8�H6;^������xwLy��}*3�'Jێ#�5:=
�����5#�Jr���+2�{�8�[���>�RWf�f\�>�uV.�X�������Y�Lc�hQdG%�U\�v�������_ۜ����Mx���_M�ҧ�y����_l���9��(�2���0jĒ�B��q�iA�.��;�7��gmC�,�!��e��������{��܆u"�v��������T��ެ��Fl weO!��g��Wߑ��X#OF� �^�G�4����p3�|�;��f:� Cw�TO52>`g�f� ^��s+�����y�hzi��k�?N��u�w�6�Sw�Ζ>�; �A%�-�x�<Y��U��vv#�C
���LuBw���(��7�[�m�M8'�w��tL-<�"V>�֌H���C�����ښ"ut3KWUB�0eCM{n�23Ȩ�TFt���� ?��I�*��]�F���F�of��"�uK��&� {�O�C��2��O�3�:=��	�	����΍��"�:+�W�_��A2@��E{TX�����7q$u�f��8�%N.�23�,�*��?��:�p+֜^�bv2ZD���	[�$lğo�n���*\�i$	,W�_��lF�0`N0���n�	S�{~��sX�(���d�P=Vv�bб�{*
�#���\T�"���<�Mz��a�"���٬o:��=�È����Dg�����oU��qN��D�@@D�*��7f���;�#����ľ�*�8m��b��fCo9���}�؏�}�oA	�� ��_/,w߅R��˚*��c�`g=&t�%�d,��"\��w����M�<���$���� ��է��jg�;J.��
�0�����2�(��r�ҽ��B3�ϣ�()W2�gQ&��y'X�U�%�Xw���+�\�R�q�7��(Â�a�C��8W���<V�sf�v�K̚�@��P�l�5��G��#������.�"��"���(؎���`���p�N7�����,W3���k��j��9}~�rn���	}$��6��8 (�B�"�X�C��v�N�zC�L	t��j���@�W�	�l8���E}�"?6���M�������o���1�D3�O��I�S���8�ם�̢B���Ip�8�c6����v4�=��=���]�.�_a[���v�O�,d��I�3�	���-���VII�PZ;ۗ��_���K����%��A��#P��Aڜ3r�f~�@8)Br��M{R�|"P�t�����li�U� ׭�s���a�q�[���'y��d��Ūs��=3N�f�1�R��0��<%���G}�r�q�����-TN��҉��`9�R����0	L���؎��E�hV�U X�]�m�|�aȭO����^[�?Ū��)Iy�:=P����P8j쯱A<!���j��	�@�����-`&�b���BW��0�:�Y�N�gAE��%��?�+�s(�n1?W�q�8�L�"�d]�q�㧓>�=]*!!��r���O��B]q�+k��?�l�����x�Z5�G��1x�k�9�^x�J��DD�©0>�<g2���͖��䑱AzpLg/��Wj ,��ڦq��	�2�BU����(:ʵ�^ؚ��Թ��I�W��$q�w0kH&��-�����GՕ��{�$�Y�2�N��L�$�y�;�a.����Ԧ��$�ŝ�|w��ٙ����q�6�?hJ���:e�IdY}$��V��
�a��;��(T[����Xϯ�0t��E��	v��R�������Y�:;����!�Qo��hqs�ϪDOk%�y v�yym�V�[E);��]q�k��n;��!��kM�]��E��h��3�N@��gh`�I���p�R���vK���2�}�Z��3�J`;$��YipJ�|��Ӡ�+��G���2s�d��.�{���3�r m|Gٻ��Ǫ,}� 3;y膧���-�5&\�Mg/N�V�Z�O��}��jIc �9�CfA��3�P
:k�/&lÀmo�m���+�7o�V"��y�B����R��b����|�����'�L�_�t���f	A]o0�������B��V8�#`�ۻ�q'�#��`ӭ��U�6��j��gf����I�m��J�C�@Xu8��/�`����z��9)�,8�0�l�z������y<���{�c��{aM}اeEafN+z�*�t�����}�Ǭ���}ґ��Et��� 4�cw;���d�$��z`u�f�����ћc�8r�e���0@k����)�-�ef�2u}��-"fkg[ K�`	�V��*񪕆�#\3�Q�Vv�����ehC�>�vTE6粝Sjv�wc��y��$.6?��+��:D�M4��L��G�] ����
;���8-��,	������xb��l��Ö���F����_��q�119���#c`!�N
�Ɣ}n�g���`�+�"���-�EÂ(bf����[^�s���E��W�~�L=�.���sN��i�P@�>�dnH�"���`��>�\z��|��R�M��y*����s��Z,ξ��n�%|�Z�$�Pķב\���&,D���&�fj�o܁�]+3P2X���Gj�Lm��ϭ�x�)ʪ�5_;�$��\����a�C���n�C6�ON!�n#�COR�][�-�
ț�B�|)i��&����6�Õ�>�c��t�&��+\�m�H�g�ĳ�xƘE��0$��\� ��G�!��	����ܓ�e��I(`�$DIz 8qˌ"�M!�(�Ku���;��_9ܴ�wz�an��a@�>�(�}����Rwę+���y��l��s��;�Њ�r|�.L�%q/p����ڥ�֡%_j4M�ph:&?F��S�2&�<�JjZ���V�HA2���	��b׼�8�����Ą�"��=ѳ���IR�� �n��g:]3�%���
��4[h��'����1���}�N�u08���G�}Z<q�F��ќ�Qj��fzE�"p�l&jU{~�B��O��'B�N��$�x[Q���
�-����|�$B��`J��*�1%���HN����C�9�$R����p�Mc��RGյN�-Vnk[.&���'�@Ϯ��9�%��6IzX�72_3��;��=�\�i�O1�M@̢?5݆���}�v�S��`�
)��gʸ�n��Γ�G�%��CiM��=�Jot��,�7;�������^qZJ��.������6Y|9*�o&�� u��m_�꿶P�L-^��V�-&�AO942�7���c[����T���E���w�o8�����8<��fS��6R���|���S��2�����l&%G����OV�+��p�H4�$��RJ�
Hs&����[M��VX<o�*9�~ � ���Gcs&��'�>�%�}��!�s�o���S�@:#�����u�s�?#��֨Ƶ?U�K�i�W��>�Mz�N�?�h��r�����F�6�1Sݮ��R� �rm�'8�N]䕤�U"p^�,:����L$��-6��f��!� Kӕ�.JD<9u�GGO�?k�2����||�Ԅ�%VӀ�p��.�ߓ�l�� <Y�L
\�LU1�Q�3�m�j�kD�a�lY�3{���Es�i��K�A�e�3����4[�u
mcb0~��Sss�M��`�է}dI�8�?���H�f�����K�ؒ�8���E^��Mn=F2:���6�4}Q`u�����, ˝P�]O�M����<��u_�=k|�c'w�,N�Z�P~�]$�r�]�ɓ�K<R�:H:gA�43�����H�_u�nr�~E�^y��"԰r�:UBD6�O�.�O���4T�W���\��֤�0���&k�����b�?�?��9<����78~� y-ކ�:�^`<�� �.��T��͵Z�op��'�,���?4�邿5�ip�v� 	M�ZdH��M�;�~�/v�p�� wW�2�l6��_e��<NT�)bQ(� a\A�rɽpY'?*U�����f��l�����V�vb��[ǖԒISf�I7����[�G�:�+���	�"�:�
�Vq��K��W"Ԏ�",�����k~Sٌ��$a�|�K5M�� �&��{�ڭ����p'1�a�Y�ql����̢��E��z�*;(W�G�y�{l���~�y����|8E�4�D�xE��5�_���=z��Eu��YD!�X�b��].���|1m��tKB3�>�B߱ZΪr(�2�g���꣊	�����b��z�0c7b���P�:y���'η���TU>yzy*�GEj��6-c��r�ӱ�(����\`es�Vg�0��|*"H΅�t�D��'2s�0x@�U�܍1�5��mEĶ�8n�kw�*�!����4�����5��2� Ү�~ �x���Sf�;��m���������8�����n��&��˓ZX,)��<+3;K����D�6���[TE���,���YyI2�I�^�97Ff��C:�Ga��/�F\E��K��J�fVr�W�n�{�q�2�s���p?�ن����.)�$�oP�JU@���@���*z�5	D�"�X��,���)��~t��f��E-s|���LǬ�9=%��fC4αo�d���O�D����ڎK:���,��d2���8�Y��X���?�N׈�X�f'��M����u�I���O��kc����C�y�M�������wi�� L#�OS� �I��=��@p������E#�Û����LY��i�P�V�z�u�dF��7�qi�Ac`?���K�f���� �{��4Tr���?Q�X�@�E�䤃2Z=WH��[�0et��)ft��h�����~�n{R�w�.)2[]lݜ9}�yaQ��J��FsWL�)�	��؄��puJ�X�V���Eqa5�^▹��C�����Ƭ�s����7iQ�ࣼ%�Ƌ�*�^)��6R�'���nF�(���n)���[|�0�"ikvN�>�f�!#���]�!M��\뽭:��-"w;l��|'�4���.��4�!Xv��G�&���{`��no�ɇ���~�װ��M��u�Q���.�⁙�DW4L]�eV�p��[��=P�]y��<"@�g`�7Ŏ�k���A_+�֜�Ͽ�4�D"��ԗa�6����(��	�l��X�h���2봗m�<-k����m�/������f��~F?����.��2��&+�8p[A蛡�����g9�d�<H�B5�w!����X�аX>�ZB��bhh~j鲸�-�f��5Ę����׮<6\��Y��q�1��2�4Z����D����
�0�g�wP1�:��=�O�}���&Z��)W���fމ6p�ҙ7-�v��O>�Y�䑏Mo�Nr�qi��ߦ���P"}�Fl��]|��@��?��Q��<XV W��]��,�wv�0���t�嘥�?ye���wV�ݢ뷒	]?.�Y��Gr��G��y�a�,�sI^"�UˎX�϶�xB˘��Lc�yC;�0�WL~��r-�CY~]�Op�ЗT+Sܴ����k���ys�v�7R���r���X�)��#�6���l)�5wď��kV�nh�����ErE��g�Z�N%��#��܌7�ߍ�m�5��u�y��t�lg�����/�����b�0�_�%)�0hX�:9l|�(����kv;�i#B�~,T�������x��^1:�tP���I5Swi T>�(ҋ2@�u�m��L	c��| �yzy���	K��wH�������Z�`|�'>+�ꯅ�)��������s�?S̈́ �$���D��5Oz�pQ��
R�<������vֹ�2͆�I �sє��rE���)E���>��Ӡʹ�����:�y�5#׿ڈ��l6�v�܀7��e6?�գvqN�U�Յ��%W#>�3!���ŏOsX���J��:;OŻ�`4�T�]��v0O����4�^�r�Q���\1x7s��<K��'n�w�����-�E.�����{�.��J����0M}�~��]zkB���+�Ճ��	Gn��l����kzb^�.�]�o�L��گ�!��T�/��+�Pѝ���3��ԗs���I�s��Ԝ{?�"�HS%v8�����vz���}���p�����^%p��a��c��~��vE���U ���3�x����z�%Ç�^ ��_Ӎg�5�K�zC�j� [v�3;nI���<Ľ�J:���E��~�� �.Vᶋ���s�d.G��ϻ@�`N��f�����UϤ�Ǵ�r��˘R������+`��R�^�=�M&�pNv�y����������@PN#E����a��\��9>��7S�����S�+.�8(�#ɓhb�Y�8�s(�t<�-u[U������"�=1�P��5� ����l�u��Ϧ�;�#�cT�`@�uM&=I�4J,������J0����ە�ͫP�Q�L�s���ժ�`H��%#��r;�2Ǖv��[kצ��!*���ֹ�-�W�2k��'ܘ|��s��0}��V��ѻ�Q�$եmlŶ0��I7��� w/$A9� gL�~���`�t?5xe ��<�ls����>�����I �[����"�����_�&K]ƽ9t�5��OT�=Q�p��ޅ밷um��V`���Z8�M��]!e��I�8�X����xw�jjũ����L���ǣ�]Z�+�8��Y`�mN�Z3��
��rg�vl���ǹ6��Dwi�uPicf�*��;�a2���d���u�{Ɍ\���s2}/�ZAH�jV_t�Q���9�r�>��]�B��$�@�h�%>��NY��ސg��P����֯C-q�0�� 1qÉ�5�y���}�<B���?g��v���F�w�73Eo�p7�y�lT'��(ŉ�
	{g�`��@�~��� e��a$<����w^�.�%�Pij�R"V�+|�~���pk�(�%]��	=J����Ph;��&�
#�ĩ���m��Bs�W%\4\ſK�h~a�<��E�\�I���e/t����<��r�I~>�aX��#)�.��s��Ã��X�6�I�u�`��9 �ԠRN��PBGn�+�u]X�����*��p�H���－��K�>��R,��x���)1���,�dv��鿖��~���#c��i���΄|\�ȼBF��y�#z���ʤ�Rt[�/��Q��G��x ��k���#D4�0���jg��D���%ZdN~ q�7��tpOk�k�^)U%eX�<#�z���O�O�kʏ��w�êi���*�o�13Y�"���'�̙CR×VK�%���'v�^"]�>֠����u��*[�(�x��������E�n|y�P�m
Ѳw��8j?;�W���Z�iw���g�.p�-���9���^}8Q�fhhi�0 �t��/	��E�Pj7�k�-�Nҩ�d�x�-�Q5�[�� ���j{� r���m5�Ƒ]��ꆏQ��.=�XgDoj"<��Qkt$F�W����w�'2`X9�Z��0)
�Po�$�HA�OR|֢�p�Q���"�_,o��m�-,s�e�}�k�k�[&&&�Ѧ�����ZL���s�������*@%���߾�+{ʴ�/���ۏ��7I�j�*�p��&��	��wC�1���#l���rݫ|Ֆ���O�5J�?�!�n뉐!����X_ ���!W]3Ϯ,j��o�!r�j�S�*i�uD_����N{ϓ�	�.���ҳ�%d�iM�{�h��Iʗ��C����3��Y�"u�N���ɜW��. ��$�=3�k��)4kqq�>�=�����nx����W��D���mC csՊ4*=Q���0� �o2.��V��Q~����1�ڪpv/�e8�a^#TS��: �NZ4�yY�sv�3Ȕ����hŋ
؟ [1MA8���¦@�h��t�	�Zߥ��$��@�~�Ν�G��\w�ѵ�e�v�@�d��g�c���DC�:��5�r�p0�4���d�-WD���~{�;Ųm�����$D��3�=g���w����xz&�|KMD�5�
g���^r�� ����G+;��$����8{�Y嘩��)�Ҽ���(�:�!�d�W~�)�J�bҺ�1?R�N�h�^�z�Z/h81��I����1����e݃��״]R�O�(P�J/H[p�p$��*�T�m����Gz�br�`\9��1���b1�DNЯ�Q����zB'��
�O|�
H��_چL�2 �C��e�S�jf����)l�=c��Lf���p���q6ԝ~�d_��KQo���u��x�b�7�5hB=�����'M�" TGpj��� �5;�'Ў�I �*�nY��x���X�/�6
�iv�4�Oy��J	ͽ��(K�7��hbp}�>Ĕ���q`����ɧ+K�֠��)��"s��l����g���T4�W�m�\��0�x�'G�c��|.*�3H�32�
�ҷ(��:0Re�����h�y�,1��s�`�3��xC����-)�e0)�6�L��>Q�8K�	;yz��Fr��B׳]ׅ�Y�{Te�3��y2�_�lU�/�>i�n�uo��EK�	�w(�p�flL�:?�S �3Xo����Ĥ2����A�ފh$�����'{m����q<���+�ɱv���B�p���w3V�����CA

���,Lg3-0.�{����f�ֳQ�.��\�y�`�b���?��`d�&������f� ��Um8���f���PX��n�c*����5�;nƂz�Ǚ��6�̏��#�Q�O���ʞ�'��G'�1�rP���V�i�#��������A!���1��	�M��3��Hx4���6��!�Q
N=���I��O`u�!o����:���N�a���3�Y*t�b�4 (�©:x���\>Y~�ɰ�PO����aO�R3`�F��	Ur"5���3���~���N���o����KP�͉fw�F�}���P��BOm?s�_����A6v�i�5i>�W��� ޭ�ϻg;οh��K�n��')(�;G[�H�-E~H�����^�2�Z�����i���H����#B�ܭV��>׭�g~�> j�L="����+<�³Z4)Ā�s�|���ݙ�z�ڽ�7�h�n�A�t�L޲T׊��l�k=�#��lD䂦��*A!�
V�/�<�.s~�h 1� ���ܷ׏d�s{Ӳ[=��g[x:e��,��ߛE���K�-�:!�o̔�o�8�����$ɗ�O�k8IҲ\��_��=5![X͵x:����e[��z)��c:zH�IV��0WdLE,Ůx(������Qn��8Z	�y�D֡�Z�r��,oz�[r����X�'��
L<d�l��Kf:��}3��I�R���.�w�y��k$��\���#pGg�j�,����"��5<n�v��j��mT.j9ؠ �4Y���S�G<��J�V�a�e&�p��QW��*l������/0Q�G��3�:^���=��� �U��~}���G���C/3�dBJ�JH������VjdKV�M��D�A�P`AK�c����+(7�}'��3�����9u#��2���sl��m�Ҙ�bGF���T��u@�<	� ��l�G�B�ѐ'�5K����q��7_��:�b��6S�š|K�������U��+����IW�*��^&y��]9ş!pq׷�C]߸N����Y���sŵ�DŁ9�gƱ��$��<`I����&K��TGI(�[�e���o�W��I>"n�����WNB¥LGQ$�J��$�������=�0T_~���1�|��:Q	�#Z�����YD��x��X�Y�e >���Jmu�6����o̗�O�A�` ����7O�a���?���Y^���ۧ�4��*R雝�
t�/���Pɏ����Qo1֪�I��<,q�U7��dev���נ���^��`"���k�kFʑ�T����Wēڵ^~����t"����F�4�1��������SW�i��R��si��t�u����c"�:�H��V2�ɲ$��On���pZ�smJ:;x,:���p�yA#�H$�4O�[OLc��9��(.�m8�5g���I��%�I��dՔ�i>�V��	�M�%��]݈��]���c�M��]�f/3#�]�RF������Lk�k��s@&�``�uM���Z����JO;u��^�\/{i�X��8��H�� gU)[\���U_1�;%��&�縓!'���>/[��ȇno�B�I8��h�R �������_�	�L��|!8��4�|Q~Xx�v�#�|��j)s(fAK8:NCstSf���ǆ]ɒ��o�ctpE�����><:���:���,������e܃;x���A�`B���Dxʭ�H���
1�j���������N���W3����nD�$�6W�Ʈ�^!+���������Y�)�J���e�oh�r�t�b�s+�X6�w̾슯��M�!	03�!�q���<������_� [��^GOІ+��(R�� �ua����?�4�,9���������F�ͭt�K��>���	Ӓl�ҭw�K0��4è��#��ڭ0^.��D�����L�I�3�j�ΘD�8V4�c/H�r�؊W���9Nx��c�׊]밝#�ӝ��s|��Z��Q���e��C�����@S�jگ���
���J[(�P��K4�����pY\�f�������!�º�����@��\��E�|d�oP�S��6�&�1ƨ�G�U�ɫ'D!�(تj@�E������\1�H���1�u%n*�s���!Sd���	���V�ĥZ��7�������;)w{��U����]��|���JT�NҲ��@X���� �EOj=X�����Wm;e-h��(��EDC���,�|u����Ҕ�V���H��cb��N��RzmO�_��<K�������"^#��(W�(�N��z�H���M���.��"=2D5�$ �
f���H$�G��K��t�Me���oq��{4�0�kx��O��v`
uuJ�"	�_�To"�op��d��s���}CA]$���}��r���Wy��q8e1�S���*9� /+5N,�׶>��y�����OwXНc܉l��P[ �tG�Yl��C�T?{*0;0#�<y����P��NNb@R��T�5퍩��4u�يea����Ż����?���f��S�OԻ	;��0�W/��)�ƕ!~����A#�`�W�~��&:��Y,iðC@�.6�9���� �� {1KN�L	ڲ��V�^�
��Z?߁i�G5L̂ޖ��!����Ͱg�٬N�G,P[�ZS��Q���C�U��e??X���H�z�g�:O�~E!�*9�-����H�APԔ"�4����G`�)�PΜ�_��G�R]ż�\;�iJ��r�5���X���e��0Ĉe�����Tp@&����!jWgY��b�o<N%3?_����J	�֢��q��#"�-���=�R��*��<�:;�)~.��@���/��{�u[�m1C<��5(	U3ܟ��z)�����ϗ�l�28�eF����E��g/���}�J]
Jc�<ת
��.c{��j`\�Խ袨~��� ?+u�5J�P�*?A���0�./ExT�v�ϕ�?T!�ڲ���w�]K�$
�:�<��D!�[��|k; 4HQ_k.!Z�Es�i)m���"W����]~\g;�q��d�6m�e��yo�6�Q����oK�azU�{�B�?�L4�.�$Tc�9�.N@mG�]���������+�E(�'x�à���n�r��\T�(=f"g�{������̴�r�V�g��dw��sf&����~��u2�6��;}8��V��6��btG-��E3�Y��zeAB���&eM8)��Xc�&��O�b��'�u� ���s���>vS��9��d�L�^F�#����U���?|_��0��-��8�2i8m)�r+�S�X[�1�v�%
�T!����!��AC~fѨ��8 k9zr���o�OR�e�_�.*��5�vg"�N͵|�w;{�DI$�t|��,����s�(m��gG�)��P�	��N)Q��A)칰��+:�/����1T>&�lZ��Z�wU���'�h-�7�*Ӱ����9_�W��Y����:-Dq�Nڜ&�lD��m>�Fe��1��X(�*+*ܾ���mx��
v�zcg@ϓ
>�9�I{;�� ��wX}��p����Ĳ��p�-����T}'b%S)be]����Y&;?���#c��N5���u>`i<;:P��#I͊p2��Lދ���=&;:�=.�fuVӁ��tod��@K���li���<P�j����Ӫ�󩩄��.��ex��'�	�x���O���q�)��V}w����BM���=�c�q3C#Ÿ��Y�C�����'-�)���
H��4����0w)Y*d`�r���0A��Q
���`����Ք����Ý
Ov����[��r���6yn�'.�AJ�L2j�٩Y����B">�8v�}]k�1�Up<G3
�"s�bb���q�M�au%F{��ڰ�][7)xp����E	dX��C��ۄ�� $͉;��=V����l����s��q0{����)||{���p��&�z��L&D�>�e���bn�4}��䫯� I�ϗ�Kj-����ϟ��5��Q��@On��^�g`귖;����6*�B5�k���;�%�odA�Q�#��+��4lw�k�}*�K�$e�ۉ&�'��ftC��xK�!J�Wg�����뱠OmğoM�LF�\�=�'[�h��K�1����:Y'�go��2��ic�i�l�!1PB�a�����)�nN�w�]:�<��R:���5��;D����/P51�"��ngi����w[.��.h�<��l"�������L@��6�1�W/:#��,����{;���|�]��Rk$�`�*�؃V�A>�L�6�ħ�p!MQ�x(}h0=�"Eَ1�x����{r=�.46�#Z�kz�e����`��:��ll�V�,����H&R�~r}����0��܄��ހ���塱��{�9FPO:{jMy����IIJ0��z5�{%}bF���.�lz��ͫQ�Q���A.ʆ	�'�b=E3B�����%5PI��Kf�8�i���D����R��[�,�;����f�y<����W�IFL��B��꣸<�_T;����BO���'R���k6�����1���έT^�)�Vr�m5�I�|��n������]��\|�͇v��2��ɛ�= ���Zq����Wq�"/��0aĠ�|X6��kS��"O�V��9�S� � _RO�;��GzN���O�[��>�� S�:�D���S�0r�����޼���Ehvǲ-�B\����g���;��(V�#(![q�G�,a�A4����ʹ�z�cZ;�9(�/���x���
,	������zt"�;^#s�N<"�󜎹�uO-����ř��?{��M��Q}�9����?����Ð���ПF��u��ge����Y4�.�6CS$�Kh¾7��8���t�:$���-�ݫ̀~�n����S�ǒm�`��Y���n4��h�Pn'�G\�u���ٗ{�r'�R�&�q��k� n2��ZW��9�aq ������w��Y=Ƃ�se&b,s��_�4���,.g������"���: `|T*����I�������i��a�>�y�d�!y֪��=��:^�	is��0���2�����RZ�SJL1�V��������*]a�"\k��ö1՟-�՞�K�!Ë&�����$y���W���_j3�M�
x���;���y��U�~�I�#�W��.5ԟ�!�?��g���Eu�`ȼ7&�4�����#�m��ar�0�\��䆃y�mDY���2��C(�lM!�]��������h��$�� �����G���;�����\����99螐�Hy=ȅ�0�D�5�9O��~#y@�=�����d����9��G�ZW^��'@�0�H�C)fe�mh`fm1���`j���)n^�����h��iȕ�E��h�r�و���(t��|h�E~�*vϣ�}����[�W4Ր� ��C�n�Y�u=��
6B�(�׉��|yg.݌8��5���pS�Ң+2uz�]B�.��LZ�K�7ڝ?jP�`�b���';�g8���F�S�1a&���*���S�a�ՙ�����D��5YR�Gb��� ��.1Ã�2�!q�ۧXg�hͯ~���6��6a��{	m/)D�;�x��l���T��QD��6�{��y����e-p�-�4B�b�+N��^����\��q{�"���b��i��Q}����^9;��@Y��d-IDo>��ښ�fD
��V�Ť�.�C���-O#�ƫ������5y�,��Hg��:7߿k�W��w���T:w ����c�5@�'i|�S�����c?Lݷl���$FȘ3��<N��(�1dU����ņ'y���L\��y�M��P�&�Ǣz��8H�q���_�l7i:A�-U7�<6�l����i��-�2��6W	�_�H6;��<�JS99���%���K����ˀe���z��r1���_ U��ʂf�l��yC�)�
���`�<2�1	���CY'u��;�2�Joj��{���O_�Ja�,hܞ	Dm��%�26�v�S5��}�\��;cI��'OIV~$oc�p�5]c�`��KCD.9WĿN�я�<��!�B��/E�Ꙇ���Yn@��2���!�P��	V:��&��a�( �I*Qi�`ɹ���9�{�L�L|#��k�}�^��ǃR�r��G�4������w��j� @U���v]�N�������ͷs���E.d����mY�s��`
u�z�w`e����߂BT1���Al�`x�َ}r��O� ��&��̭R�5�$�������Ҡ�S`�|�'E��8.L�pm��TZ6�HA�H�!L�C)։eV�:�VA�a���WdHe�َ,e����p��;F*�*�Y�B�îo�O*��6����Нy=3?P��➯�|����d�/������i�O�,������q5m";�gI���̺|�-'$GϢ�����֟�.+Q^���r�B�>�(o�=U�`�������r��[?�A��4[�^랔��f�u}#Co@��^���H�┝n�+���{��j�?X��p�fc`>&��y������>��w	��2�=N�F�j g�F�2`Q�j����rj!Aׯ����m~㓋�u���eٞ�區u�7lD0iIԳ���_<@	���'�x�� ���c�I�
��� �U������ገN�����Qץ�޹y���E�z�� ��}�z�_U�.��.^ZZP�?I5/!hT�H��!�D^?�饼�IP�t��35\�i�Jڪ`_�� ����}���,	�9�s�f&��j�xoŵ��M'G���.ʥ��=��<�f4C��䞕��?Z��o8{��zIx�^'��Ԍ�I�Qc��&+��0|�(�·�\ns3����Q2��ocY���0�&��� �K��y�:�J�C˻w�]}ex�A����Ք���@h�ז�$]�0+�M�Y�(�I�9��$@�X\�dXI�Ɨ�{ph���:�G��~�*�kZG��ن���,�/{yٚ��%(Ħ:W��f�(	�����W��_�翀:c���,m� �OvJ��;�y#Uú�_����ʁ�Xʤ*j_Vp��Y�U�N��.�3��K��oOj��[�bd���'Qu_��z��{p�����	��D4H!	�b�9�$Q��������$�3�X ��Wk�P�������[]����C�9��<H�b�a��ir,��e�/98��h>{)�v�p!��"�^�����Z(�nX]{��ݙ��L� ��u�~����#����-iu`��Q�I�k>&!Z%��B�u�A<Y���9c~
��$>m�����/n������҂B�U����Ә�v"�BXC���R�������ߑp��W�����`�
������e؆4���G�b����Yt����>ݾMc
j��r��FEI��-�k@����qF^'�!���	R���G(������ٻr,l�>���yI蚈|��.�O�:Ah���J-�mфH��:D.���6��r�� 6z*&R�x��O�ܣ���MZ�Aק�fɀ���w��4�-g)C��I	~��FК6>+�l��?��"�M��C�qDV�i�_�=6=>��a�(�'�ش���l��Ҽ�|9us�J��Y��4����a���	F\5K	_ח�$��*K�7"��f����L&
 �����h՝�(�7���[w��L�mI9ɳ'�}���sn_֌U�s�RPb�c����[�|5L��e���׼r���d�N���%堃����U�\Q4{��
y190��ÿ���0��&��0�i�Ì��c��ro�c֐	�s�fؒW1���d�e�h�)�s��nCG��#������krU%&���E/��+��i��1�%=!�K�+�Vއ��7#�`�;�ˁ��t[�����W/�E5��Ga*<�����C<�n)"��Ԋ]%��E6WW~mh}���V;a)΢�w�<:�mmf2e�<�͠B�}G�}1�\����P�s�X�c'��3Y>\��\
j%*:���|S���y��1��Q��h��Բ�.����u�:�X��&?LE���c��z�u��JbO��/HJ����U:M�l�TDk��5JCN%d-�xإ���	t��Ȕ��C��ȡ�h����t�*���~z���G+������Ka~�;<d0����l��簠41-�wOT�!���Q�2�1�P g
{�.�(g~��]�D$�S��&��k�/��B`��7���� �
��_������Z�I�+��^U�.�6DT͵*g5wߠ��4�aX���DRZ[_}͒�pVP�@6��#��:T'�J�+x��J�����^o!v�._��z	�¬n�����/ReK�0�����Pi�2z�5�vn|����MV������|�~�Cꀨ:�aM�oL��V?��t����G<�DWӾ�Ј�c��k��-rL�e
5�`�����3tv��{N��=?�]��0�W�#�u�+_Ps����#�X��@�>!��E�n�u�1 ��7�S�6������{��2!�����t�]=x�k��<���S�(�U`�&��7��WKZ�wUL�Ѯ߸*=fr\�[CV�&=)�"�" k�Vr�5L�r�XO�+PMq��]3Y/{R�˙�� g��r���*���3p�2$��e\v_���G�%))@���}CT�h�h/���'��Z�7�ZQQ̯����W���n���Y�f��6���Uh]�9,C�ʭ��r�� ��oc�g���:M�(�?�,�q�������]Z�~X��)7X#*���V�>Z��P�?\���.�+M8X�?^��8!��s��3JK3N�*;Ԅ�>��M^�W�I�q�^�,/�e �UP'P&�+B���_�UP�-T�L0�q.�'��1�B?Q�w���J4�CǹJ��7�K'/=�ƸѬc��>��)�o�n,{����+
��4T���-�A��x|�-�ڻb ^r"�K]�!�ŲA��W�~�r��v�
x)m�B鯯)�C�eԉw[Z^2�5��������
kiX���;��3��l'��`Z��kE{����}"^�oL$�pz��&|���8{sf�#�G+��p��H߷O/��D]LӗC[���7Y�����>J4����Di������q.���C��u�����;;�9�1ԗ^���_�
���y��ދ������3�e�T�(���.x�R���H6���7����@�;2�;+�#"�L��C�m�1��;�����Zo`Fv��N�_�:�0֎��K��
�k��߾(��~��."�G�v�&����1v>Cj,)u����T ߘ�8)N��`;,*����Ǝr��ki����Gw��
=`{ӷ^Qu�2�܃yB�6[�)�Rf����^V�-^��fݽW���Lh:9������w�[�=��1z��kd��w��[O�?u#vsb�C}Ɉ��v@������#;�H��P\A̷�GT�Ξ�f0��������t����(�&���Hh�)^B���C����M�2�������������&%���8�?<����àJ��n�jW�����n�w��ſJ�\�W̡�K-'�{L�$�R\6[̓��ܢ4��B6<A�9 �fO%ޢ���I8��u����KW�gz_`��aԀ'�a��lb|/��|4�Kr�B�V� 3>�5�.���Jf��Ih�X�q�����Ʊφ����� d���h�!��)�8���qjq�����%�_T�n�+>�o���܂�~R�(�Syd��s)L%���2/�#(��OH��Y�tv��c�1T����T�f�T.�s����E��]Y�
^���^�܃!�iOfH�P���lj��{�c���:�/7x4i fr����f�A�15<7~���嘡<����t+�w:�۝��<��̶#7�d�
�.�;����5\ȏ�\�����ۿ��x����?��g�K���<�X|`�X!5� ���Nebւ�.��>L�eО��<����M���gs$�ۘ�GAyεe�͠q������ix���90�t���%�~_�֞}�wœ�4uB���4�1��N�#*Wr㣹��}���/NtD��j�h�O|������&����`դ�
;�߬��bn�]��8-�"a�a%�m��9U�4+��lƏ���U�8Pgg�"|������XQ.��t��Y���[б-<����� �UMm�U���z��[Dγ��
WU�J}��^q����;{�4�ris�g�[�����Y�tlW���h0��ߪ��L��� *0S�-���t�WBL)ۉCw��A aY�I���~��ܢ���A}
��T��PB��GF�t�� \�4]��.W����k�)\+���.�\7�=�q�������^�d���t*nr���͇()}r.�'r���;1'dO�	wf��l��	f`���O=�>E��u�=�]���;�+o�s�䷘�6r�˸���f	�N����Ո&��)�8���8$tJ�P)�\�UPÁ��me=�����_|�Q�~�'06&�LВ�a�F�kjZ�M�׊�>P`�[��_ܪL�\�\ �~T
8�;��X�h.�n���&�q��I����GC������<�*�x-�<�S��$�gy߲>^��B��71!�S�[�F&��J���0�,j�!��������%XST��ԗY�m B�B�q��L��B�g3�ñ�PAu�'�T�:�i<7�$(\�o�TGa�������8��}��R{d�l-q@HR"xw����끓R�i��l�s��ٯ���ϱ N�{w�r��`^Wr�f�� ?���b�:͂��G������p�DF�~G��j�Fn�C�|�b#/��C��e�bv��S��襁��`#�%Vn�D���gn�s�ݣ��mZC�%|�;���eVvň�S�ZԈ)O��Tɚx����U�o�R�3�EE='t�xs�S����ݒ}k�W$=�����ptӌ�'	��2S�׀G�>���!L�� ��k��Rn��4�~U����]]��i��ق��C{ͣ/�Q�u�W�1����ssQ�=�$�7�X�:��|�
�r������S����J{_+d��~A�1�ޤi�gF�`�� b�m���S4��޺�� }!��x�Ox-���k���s}W����0}I�lܰ�"�Z;Ff4�a�]*�cϴ��iM�P�	B�_�wp�Ŋ�d��Z�	�!BP�H62�ʌ��yv �G�f'S�hZ���p$A�&�r$w�o]J*+�yp����\I����tv��?uH*��D	���:�D���=��0�.Mz�r�c��Ӎ�O�u\{������8r]@�ԑX���d�9z�,^QP,M���k��2���JC@P��|\����s����f�K[�H����{�!#����ǩ�=�	QMq�q�B46k�h���=� ���@���j�S��r�Iv�(�2��%r���W����4q��o��Nr���T�v� ��i�lU�{�˭�K>����7��Xw>xb���;���4Eu��F;�5٤�;����s�;��4v����bEۋL���z��½TU���j�M��9�����7���`,B�����`h����^)4U;�Q��8�t:/���cUq�����
$�7&]m���hj.sZ��1 V��My����0o�0`n�1��o�)�����h� y '�����?R�c��V+K4�L�X'�jj���#t ��A�X�}B[ĕg�?��E��g),MoEx�d�V�02@�����dodr-�19�(���s��Qx�
 ˆ��b�EF��|������Cg@���5��~̱���
t6Ɲ���5���>ܩ���,&q�f��C�z�@��x���|�ȩ�ا�1����h��"F4vE�A%���PF�����6�`H꾓Fv�BV��#-�1��{�L[��3=�nYW+fsl�ђ<�M髙m,<��bZ���}JT0���ܳ�8��e\T�9�3�f���Н�fx`8�vظ*�}u���L83���V���i�!A�B����V���ƿ)�),���v{A/"dw%������}�+����5��4)�_�b�u�.�*
X�m����E����O�j��d�Hn��Lřht��9I|͂����
�n\���X�>nE+��vH�ZlJ5�6F+�ց�/c@�{Rn�����j$�|k�$�a0\��n8k@�R9��j�I/�Z���.P]/S�\�(O������/��7����]KS��&��S	x��zh�h73Fc`�ʩ�(��,	,*E�t�-�Z^;�45e��A�8�RU�G�{	�a��O9zh|F�1�ɘ���cvC�5'�#i�w
5d<����>���ܶ����1�:��|]�ҍ��,;`ZD��5����Q�B2g1�`� �y:({�`l�i��\��,�����_-*o�y�����:l�ڵ�60��ú�����np�S?�%�u�-Z������0:f"���s����X�1��"�.��byH]0(-���f8sʓŨa�������r{��<!e��a��Ѹa������_]$��7���K9�����ʷ�_�
�J��QˀޯЌ�ފL؏��3'�)��Y@.x_�Fe��E��b��bN�<���R@E���Ҿ~E�O��W"S%�CO��c&���8����ЦTi��f��YfSo��V�I]�?���V��Šл^�s�C�9��k��?�M{�Yt鏺��P�>�
�@���$�բ�4�D�kV�&�4U=4�ߋk�y�\<�9�3�fзF�r�n`�b��,����81g^յ��!Y!; i�T�t� |�L	����)�;D#Y�î�p�+���1G@�R�����>8�{�JA�оB{7�h��Y�2�U�Ж6�ztѳ�8�܆�oW5�� ��a���~�\���� �&���K��)�^���� ��G8�I�v��|��ن���dC�C���p$��F��a�DŉF�M���!�Ow�::<��f�S��*�Ppv�.<�j��W�1Ρ���PG�~�_�U���:�%+6�%âO�p�Fb�8��9���óa�姻˾�}e|��`�H�EG��5lR�ZU�_�N�-�:n�r*��br��s@ܷ�яr��XJ��G�P�p�ِ��3@��LH��A�%��و�M�I
�.%�l�C�SL�Y��hu�T�;��
"J����ăUapW��<B;ǗN�-�/����Ӟd��f��<��5�Dx�6SY��6�}lLI6e�ȕ[l>�x޴��:3
Kr����掩T�|C��h;�e����;�υ���x�P���4N�{�������tJ���X� ~`��2�:M�����:��wo�`/ў���,�_9�:�b�NJ�ƚ�\�sG�,G?�`�B�
Vȶ˥�lw�����H5ґ��>ߢez�s��Y�Z�6tm)g4�
^s'	��ޔ�^��mZ�(Ģ򊳂���	����Yܺ��V "�AHk�2*L�gJ����������5���G�M�z���,��>6Y0�if�����
��H��䒦�?b&)b�,���[�\��'П��I}*D��-�k9|Rȓ�"-�����諙;ΥY�}䞦�]��H*8�XE�"�]h\�0����'�0ʝ޵��g��Ū��R�Јcj�b.��à+��u��jx��c��I����~!��'���΅�N��S|��7�^*'������6��j�ܔ�1R'k�Z<s�h5I�hVK����7��|��s�T�|V�e(N$/�o͍�[��i.]��׌�z���9�֘�<|mj�x��H���	���	{�A�)h������@�F$Vp�|(���4'��,M ���^���qy5n�	7�Bؼ�NVXΟC�M��l�+�Ρd����_>���utb����Y��F6�#�f�����CRA��t�j�ʧ��A}Yq�0D���Y9:��<nE��׾�w�u���ҢKt,�������uݹo߱�h�]����#�e�ޚ�������gRKc�8[� �Pg����Yy��ոb������?��f�����"��5P����Q-�� ���?�VoBC��؄s �8�x�e5�W��4پ�@4Kg�$���c�@ ��a�0Q�+Q�7!�0s�ڠ�G�,�#V��G��ۜ����T�������NY��;�tM����%�ܸ$5������Ktkz��H��(����f]� ��'���%a�]��5���]�I'�_^R�+�ޛ�
�Fil�LߙN�#ûm #�ق�:i[�@Q<�E_h;E�پ���\P�,�N�`���+�'^��w���:[�nO��H�������	�RL��G�@�)�B�9N̍��<�V+�L@<4P�ͱ@�V1���6A�f��BV0�fۄ�?���@j�\�{E�#�KN�W�;��l�U�T�g,���(^ւ�3�`o��xZ� Fs ɱ�Ͷ�0�N�#�8{OB�E&3�N[��bd���$���1��or�<���Z���N��)�A�1ֈ/��h'��|�*ӄ��K�}���a�	��Oĝͻ���~�P�tt����'!��1���W���+��&�{viڟ0����.��f�+Dc�?�j�ˏ/K鈆V@_����Q��8^�F=�`VA��wR$��v2�j�2HЭ�L��>�).udTm�� �5O�'"2*�se�bW+>s|��Ot�$k҃� r���y�ы�UD�Q,��xXk,V9��U�V���]��i�(�}aܢ]ּ���羸;2E*ON�"��M/1Ĳv�gF-\��~�����V�/%7�G�P4���pa�9pޝ�j<�R��Ԓw�W>':��#�B����a�/N�%s.�s���P�H�k#E�'�����5��}��IU)��?�Z_`A�S�/  w;�ӗ�k�d��ѽ�xN���t�:?�3�k��"�[�p����Epo��zMր�VBx���9���H����K�9�"k���E{��Ƹ���U:��e%M�Hwl�A�ƍ����h0���	P�K��ܢCƳo�VbC
����gZ���	dF4w�?KQ�,�v��4���S�c0{���[n����)�D����6�u�o`mO'}	�5�,D´~�&tH�YC^�	i�+q_ldY&d+�����?��-̀�}�o�69Ph���0����(Y%^�*�K]��S׵�-�mC}[�m�¸{�ͺ%�S*��P��L$����f�l�����>�y��n�/8g��a��<]�&�9Q_�t��tIn?Xn�æ�Gʉۿ��Y��T{�g*42s%A�/�c�a��NĆ�a�M�n�d��ԗ�6�J���v�lm�R�f�U3�.x���S7%����@^[��Y��Kē�ڌL�!�u��Uw���Wu�]��'=����`X��A��6̤�
s]��!�P� � Tg�W�z#�5�]�5�4�L��8	�,���ص0�r�_��>�=1x��	�W��2bL�(�N�ό���۱��0�����:�<d�O��f\��Å��f�cX3��T��In�މމ_+�>*q���&���Y�w�O�����9'41���y�Qs&[\�3%kγ�(ȯ�687�{E��)�3�����빌������[z���,��2��IH�J�^���s��G�.r�>�;N��a��(/-�J���J�E������_�B����J��R��5������i2k*&3���A�xܫP��_���r;��1���eg������'�ԒU�p�X*���g�{�Ȑi��\�~�Y0���;��d�u�%I��A���Tu7)'J�L��.�!���Wa��
[���exHZ�������<Z"*���mt�ME�.������bWc��cl��>(�گ>oG[l��f�ɗ�����R��+YY�?n�'P0	����e�h2������^�<D�V��w����Zuu]���;�H���BLMte�<�[t���)���-^��x� ��d�6�1�h�S��h$�"�Zq<�����*wq��+L���Ld�Y���T/�s|�^]*����!h�'"+{��J��~��^�Z��ܠ�du
��#O��R
�!dM�3��{C���<��n��P�{ͫL(=��p�Q����*'YZ���(b��{!@�gU�&�.F�8��o�ט� l>��O<ڝ�Uf8{�oEh�E������<͐i+�<x��fp�Yؘ1��k�eo�sFM �DE�[-�bI�]b>��B��k���q�\|v��Eg�#�ߠq��5�ڧ�UC�MX��wNtB0�?f�������B����E�r<,WWα
��r�D:�z�{n��3h��������~��-�q�I�?F�H���/Z&7���D�;~: ������4�S��܍bQ�Ӆ>�����)��؊����1r��C9�i��vy*����yN5�.��v�G �����V�����>h�������.�B�U� �^�w��C��~�C�T��%�zYe��6���EA�E(]>�á�ۙЮ��yL��li�m�bB��%,WC;T��:�.
7r;QE=�C!)���/��/�m���!��� ,����&���~��^��2
>�	����I��qB���=L�G�K�KV�؆��UH���`��@��e�J��6Naءp|�焖Π�Gĺª3:'[�Q;��[[m;�j`ӯ�J�ry ����*����]�V�(���zP�9!�D_n4��������z�0h\�hG�y}tAx��X�7�F?�����f���q�[�a-6ܥ����!0
t���p�A����R��[oE���I ȯ����hw��!�`�С���ή����$pطA�OM��Z�Uc�����R`��Ni7]8
��R��I��dJ
� h%��i�n���)p�ϱ?��mTwa�|]P�f7��g������bU���y�������{B�هykF\k0_V��3"�M��G�	�pɽ��ն�f�����\�57�'�Pȗ�;6���Ok�ᥚ���Li���W97UBD�V@h�|;�h�B�E��.]���h�0���D-6�N	�S|��:�3�@���zIp���ud'��8����rb9Z=9-��`�|z,�˦�Ω�i��|C�6��!���"-�GR�KA̦�yX�
 Zf�.��e�"�I>JN���7�C�O�	������k��V\)��I\[F#�
���#�������^�_L��A�*�7M�3!y-�x��e�ֿ�i��t��:ȓ���~%���V%�����ªJ8��Y��.*I�`�Y���_�^y�A>p��\h[c�LBZL89c&B����_Vb��'��ϭ��r��D�*@��n�iփI8xoX�/�j!�ʟ�Eh��+�]����l�mZJA��e��c�E��vt�s�O��5�P�֏�$��8M!0x٬L'ž=W��Ɏ���Ď@�@� �ԙ=$)_]{]��Ew �����=��+,�h���oF��e)x���K0!��WwcY�sE�H���h�^�\����t��{����Qʒ��>+� =W���>�r��B����
0��C��Iyy���5�gi���.����R��_t�bN�trKY�C���&/�^�{	�״��j� �_ܚ�fA���^-к���v��Tey�-�g��Q��"�������w�'.(-,'~��J�~�rD�� :'˩/���®�߭�N�����kc9ϣ`�<��JH�]��������B���5HJl�h�7�������<��k��)pT9�f´�-�Fі�Q&�{"�d��uLp��̫J��k��":��W$
S�SJV��O���~�A�p�?�8�U��(T�z.DK��ʕ5+�^�;K�80u;�^�+n�O\Q_�]������h�߸D-�\�]6�T�p�lT�eg�ا�q Ǣ���.v=O�C��v�c^�<_jń�b`�+���_�M��ޔz>"��Sy�g�����-1��V�o1���M�S	9�?�u�zq(\y�f/"�+��c.����K,�������03S�㉅%�ˑp ��W��̨�Y����{�M�t��4��ݦ|@nn:�1�@͕�?
�2L��I�69�3�O��N�/�w�m���V�ʵ{�P��&{;uYscWx�5'���}�/$,�N}֧�����o��,��0�E)�ҵ�Y��>$�����+�&f���!�4���T(�w{\x�Oxɂ�����U<�|?BG�fԑ�s�t����ݥ1-Xl��j%��WG�8�=f�]��D�w�h����jh�G6kD��J#��a�-��n�׎8-��%4Rv�a��S��M�\�Ng��-�'~�dy��:C��	ӓ�'��ܗ [��-`����������:`���׶��������[�3���OMU�U��x�0��C����q�a��|Sf{=}@���f]�QA��ф����u9a2Ó�ش�5�Oy-�6�I
�L�"Z��S���&�4�1j7��<�<�_�R; po-m�|��{�x�U���j ���#�-����Pv��u��螽#����i_�����7����/�c�R~N��P�"^u7g���}k�2b#J�yG �Ĵ�bY��A̔\����r�H����A�Ѫ��Rb��y�&n�jF5VD�C�tn��L�C�H�d����<q�E�=��=))D��+�hj�.��bp'ZX��bi�R'�~D�f�ً��F�2})m�<A��x�B$~�č!��V�UVO��i׷/���%)�2!��tާ)'����Y�"�cC(Ȅ��E�'rꛔ6��`k�Į��t�l�K򚷼i�|Bk������4Wx}O��	Y�z~��f� �)���w�:qI��B��b ���N�Rӭ.cV���L:�J�PuK��4�8�~Yc\R����4�~&O��Zv���xա�A�qP�Um�2i&!�8\ؽg�� ���)W��6	F(-%ѵ���-ʶ�O'āt��3�G+�Dc	< kt�����u樏o�,FT�u#�mm��d)��/�joq�}Y7A`�����>j[S! �GVB�����+r_�8��T|��uÒ�G4M����<	"u����0h�R釀0s�
������|�`�p�J6�����%�SƎ��=Lh�UY�g$�&��_��A�
5�[N�W@̀(%��~/2���I(�6�c�������-���SgrF"'��)p���NC�U-)���c���l�ClV���"�QP�FԠ4��ߦ� �B(o�������"�YŉA��ȝ��<0�Ϡ�IK�WexKy}*v
ew���(*:s5,��F8�
uܳ�9zȑ"e�����xi�B�x���<a���M{�Z��v9�B	��a��;[��@��:�v2_�1��j6acD���0������J��x���9���3�A��n���q��s��_J������)�z`f#@ԫy *���0ԙ6�ݑ���Ϙ��̷Bf����Կ�� �V��Ĵ�nW8�ӑxLAKv�?$����ñ�>F�㐧b.b_���CI�8�u���gw>�"���ۅ�'vQ����8�UcH�V�l%¹������+�A�:�׆�;K�Ç�L�-)�����'��h�/�M���T�-F����9�8�"�����sZ�������09Q��+�r���>�F�A��#���?Ĉd1�I�<�rJev���oIЪ�KДN5��w|���>�˯�'+y5N�bH%�;�Aߧ�%,<�7�B��Y��&�>�Lbc{Jre�U����X^=�pRg��Z�a5ɒ�p��4�����F�X!�*���w�{���J~,�G4#��{�j@�����nI����Z�6kN5��-  �^[�:�����!�|R#A̪��G^q�E��դK�ήm5���>�-˾|s��aQqλ1r������	iE�ŲH�d` ���|q�aq��66:�k&!q�A���C󲿑�l͛�7���p.u1�+�Τי��9�N�d%�ȇn%��ǆ=J� ��@���kT4���Go��:�^�cm �Q�5��"�e�L�)`ɻ�)%���:b��XD�WQS�?��k[�NcK'�g�{�p�5���#��8��Z����Ka�����IﱗJ����sZ>m�qـ&Q���Ј�j�C����vjO���Ν{�f�j�p��S2b���^��>;A�s
���S #�QQ�z�R�5��C&`1ޒ�p�]6b�ʑf�jgq�k��M/FX[!�ׄ7��z�ޱ��v��F�󩩩L1���F�{���>�r�V(�,����>�b�����,b\�.J��.Ik���`�)m�'�h[�r��÷�S���tv:~'.G��E�:�:�&����*�i��~��W`�����^�����zw����V�-{��8�8�����m�����1��3'㏿H���`vW"n���)�5�����g�:�}�0�.VB�v�NU/�~��A �:˱�٠�h[�LLt$ԗvu,�9��z���vo�!WP�n'WG-<��"FҀ�!�i�ݛwm���Z� �T���է��>ٓ�/"�(��9�T�v�ug������N/��	_�"An?l�� A��w
���[k��#�-�ʨvI���ۂT6�-3�_��Q|*H3�ĕ\��47ds
��O�U�Cw�M������[w��U���G���z�>H��������CC��Ac?j�	³](y~@�ǯBs��{8r7�Z�{��t��^�w]PV��vѕo�[͏���A$��^�����Y~c߀��߄F;K��������`D��\ÕFX�vޘK�q��X��B(	3��W�ڲSɢ[�nn����A���U*��!�Pp�@ɠ��(!�-�t��PKϪݓo�PX�]�����i���FI�Q�����*FHnD�����땚ɯ����ͽF MG��#؏�alי�#uÃ�!�V
<s��*�� 
+������i/�_���W�$�������&��pU���#��0�i2|��Z�; `N%Jp�$����9��t�d��#K��3���f �nK���08E2�i|�=�sZjj8a0Кh	��|���E�"�W�,1��.�O���B�
kI�����c���YS�j}���`��C���k��A%1�y�d�?�G?Zjg���4�w�M����2:/�ᐨ{�&�d���9�I����;!I�v\����+�,��h WH), eyC�>�6j|�@Ř������� �<�hn=��Yia,o[Ԫ�8!���5��y2%v�\s�M:.6��pvt�I2���� �|�:ぉ�&ף�@�L�&���Hm�T�x*+x�|ɒ�V�����S�PUL�2�U�)��֍���b�ί�_�E1&SD���.������ցd_��!�*���*��?̅�c��-M8��栗O�]�=���C�B[F:-h`GF�̋���kT=��εoц�	�O���|�V�~����{b^�H-6M46<z��Q����/�i�����Y���%��nʕ;�gL�8�3��w/�.�Ϋ��a����/{9�i�u
vIY&�)
ާ�4n;LM�~�N��<�joXjH����>��{�$ۨ��Ԑ�h���r|QB���e�hU�#-]�h��,�)�D)��S�]�X:<��l��K̟B��eȟ��9��_��%J2NVn�؛3��O��a�H_���&�EwɝG6�vʬd��#;��R�1�E��s�q�u	�a90��ȳ�y۲RP��v�v���`q������z�� _�[8��?㣗.���_�H0<+�0Fg&!��eof���޼'�����N�bKa�2�dq�~h3�f��`��Z�Wb�����8n�pw�Τ��^;��+k����:�;p���o�dHFt�c��c� �Qkd1U���[�ݩ����l���t\���%z�Q�c��s8����9E�T���Sjڈ��z��U���ʹ�pM6)�<�_����p�M��p*#Z@O+���K��a�\�k���P���vc����p���S���TU?�\]/	��[b'��_'7�]>�f%6�b��f�����fLL���o5aݳ�R���)�e7�q���k򸮁�O#8��x.	�'���2���>=+�s�剔C��0��W��+�������$�\g�<b9���ƚ���4Kn�=U������]��Y@8����+a2���v�,Rں�I�[���� )�.�q�S�0*Vhg������f��驶�p��J�K�r\�m�MPSt�و�s�0�,�.�:��!C�]�5b�_�9�RV�� @�;�H)!�.i�*H#$��u�G��ɖ
��Ξ/c	j�&������8"m(�Y���iC5ٔ��*s���<[�, �)M*�{]Gch�Y�&.C�8S�PW�/�ꏱh�Ħՠ�4y,��GǕ�P��~��w���7��5�vE�>fm���r{����M%��_�ٌ��鬻��po����P!~gl�G��9oJ"ϥ+0V'�z���H/��pXO�x(���4/?�& �|(y4����,]���X�F�l9c���V{��R�A�é�ū>jdI7?�ɔ:β��.�B�A�,������-I�uDC`��0��k�d�p�'�{5f�Խ�R����h�1<x��L[���5�^��<qU s$�6�e$H����xrݳ��w��Ć3�� mV��� v�j��C�/x�!}�T�Zn	�|�>Ʊ�[���R^�M�!�x��g�(w�p)��ڮ�<A{-���Y؛hF6QN�H?�:�
U(_OF�oU�o����'F�,qJ[d�P ӟ*��R����0Z��IE|�n �O��T�����Wܹ�K!6V?B���	g�wN��qJ�����a���k�t����U$f�[�=��n&^
8�Sv7SY<��� $��Ì�8�/�g+�ηX�Tz�[���v>!T@�ǌ[�_��T�i��Q�!i��I����}�gҼ��k��-��F�5PE�2W�ֈ �몪$�s�i\�M勂�8��Eb��6�b/R34�@Zp~���z��%H�v�"�#`-�����@`�-=����j�z�UW�}؈���ڠ.�����f�R|Y.� ����Y�h]�P��B󗚙�^ ���w3|�)��k+�Y.�P�M4�
B�MR����&O���2�l����I�y!���������B"�~�d|ڌK���kG���	!�1����Q[|N�b��xҎ��,Z�-�R�	>T�1E%�^8.R�-/j���@�q�5\�OI�U��?G����0��p��u�[Z:D���=��KF�e�>$���:U!�B#o�AP,r�4��f?9��y ��:t΄�����E����k�gJ�M
�������S�.��;F,̝uSG _�D���+JX){�P�1Ʀ�r�}ʬ}�d������_9��ѥ��)9�j����K<��R8-��Ŵ{�$6�K�����/`�M�Ρ��Q�bBt����{�7�iS�2�I:Ȟ�l����kJ���^���8��R�1\۽�Z�9Y)tK!�ځ����顥fʸ����BYp,����n��&�����P9�>�KĜ7Y�֍��2��#FP5 v7٭7KAb~�(v�B´�3M���	sxɲW��˲ؘh+�Lk�-����a;^ݹ�^.��XlQ��A���_Mݬz5V�e�Y��}��dܒ�.���enT�� �%y�+�RhM]h��N �`�h�L����ܤ�d� ��n�7$������b��9_��Z�T툋�(��æ؂�T�����	�o#S�b�Ư�����oR��ut�m &�,��$�z�|��&Oe�I�+��:m:V���u{�K� ް}�)\�gp_�;�O�4�r{�8�h�f>9�x��"�Q���ץ���aߕm���
�r��;lL�~t<�	q�b��4{�|`i��}�W))��XV�S:^̪x�NS����0��.$5�q�N�^{�!Xڷ��E�������V�{Iǰn�Lѧ~������͠��P�χ������)䈗�����4pp>��1���dc'���mﻣ���-�����}�kE��N���@��4m�C�.*D�^��n�Ԡ�u�*ULZ�Ƽ���b1��9
���4?��ﻋ�yf�^��=g.���Jl_�Q���,����P8�?7���ȓ��q�b��*��oc���
�a�����II8��œ�(�;d	Ʌ�qlEm/�e���R�C�]�{FI`��� �U��OO���ت8�X�ҙ��)!�v�Y��疒ޞ�s�L^�w[$ ��̰Q|�^�y���(�qTe�[�+��:P�[� Â�#��r����@I�djU8R�H�/P�Zy{yJ�G�.c�.Ζy10̾�bNכ�k�w�������W_���"~A''�-�����Q�{3"��y B�.�x�^�SS>EΨ������Ϩ7��s�6�����SDמ�}�w�Pg?�Q���ރcG�#��6������9쑛�]�J�x>��z����+��`�z�>S�cntw#}0���pI I#�2�:U9Į`�k�/����Yk�
ȁQn��ctr�n��5X�sC2-m�s}ؕ�M�<�X`5V��'Es���q�NQ���P�͈5�R�@�tBG�\��(g���)�m߬�E�l�Cf�S�@�I՝i.XA�9��Ѓ|���ߎ'����_M6��+c�(�|,��}��m14�X�gs�My����WF\ttEU� �T<t������x���@��Fx#�\�f{�S�p�ȩgQ��ک
�B���˔�qfhG���-?8#����	�:�K�݄��!�1
$����N�A�L�Ag\��j��=�����|�2��T���ݿg%�:��rD�w��0;L��v���L���}>cÝx��&�4G��G�d�-�H4�;]��z�����R��UX�CXߩ	�R�64�&&����Qc������Q`��eh�q$�	�%���i}��M���h0�� @o�����5�5݊�v�(Ħ�LP���Z���\��{��o[���N ��'A!���C8�(�#�����!�<�j%��Y�И%�$h�I���IU�K�/�֓f7˕q���ox['��ДzV������`z�ꮕP$Mc�4�-�N�n�%����Wa���W�7d)%`�>=S�����AA�L��24�3�Í@��,��k���f������g�����b��0��֊&�8к���*r�5J:�I��U{G�'Yj�9�T!�ש�U��rio<�D�t@x��7��;��j�'h����i\�Z�p��s�1��Q�7�v���Kq�hFԡ戔��P��+�K���X�D���7/ɕ�G�a��Y
b�Τ�?s���O����]�A�������#����51��.:f���қ}�r�-_^�7�ΕC9T�!z���H�\��������z�S���c� 0�z=��x��I#�������dY+�pk����K�ۻA���2�������vT���W.��we�-a3p�ˇ���&��:w~ʆn�z�=e���TZt+	8~�u"]�m�'Y�N�}L���|��*�Α��+��=��@ ��Y3i���}W4�>]S����&su|��J#fO�|;���sn�v������!�@�k����|�>5�0�{"b��ꑯ�E���q�ߞg1�)��9�AB�լ�����:OĠ��P2O۟�B�qa@>�`�m��*{�|�m�S�~h������a	A�P�K[)�����oՠ�'��'#�ےkI�c��D�!Y��U�Gla@@���e�s[gAt�L]X��L�#�c���^.{'<�	TG�'쐁:��y��8GDS�����#�
�������YJ��Pftʡ�0��En]Ľ��i
)�t�`���m�j�UA���L��rN�H�f��ޗM}���J+�{�h/¢d�M�T闎��vz���D̾���HE��Ee��k�d}�4�O�`�z�H.$k�m�ח�վ���>��� s�
�%��vCWF����ߌ [���.�[��5�f�2A9.y�s��2��������܍v�s�ӅR�c��d�͐�L���s(:mP�&��+�G��s;�v���$�i�F�.D�8\�2�ʩg��_7�q �p���Gzrі�g�	��}���u[5&Y/;XJ� ������e��r5M�ي�+d�v]�/���(U��� �+�����])*���\�me�?��!��r���]���a��3.f­-���<��Z��Ti�E<�y)�2�F)��­g�tӠRz�6�ɚ��촪4�<m8���'ۑ\;�
���lfq����: k�4tv���aҰI����O��wH4XrP^A(���U�0�%�̫�yY�v5��|�$��������N(�uI��л�����%-�{f)��w����)�;�!~��1�"���H����+�@	��E�(��,����N���vBAKޞ������E�m:c�_�!��4)��Q�bֽ��E齣�M?u�y�+@���<v����thT�R���U��D�P��1,kM��79��jR㿦�VSn#l�31�s]Y[kp�ȡMY��t�9���7��੻=�|W�V�<hf�#W���q�AXc��îr �r�x����
 �� �v{�ja��(�����HP'��#��Um�V��8��b������n �p!����,���"�2r� ʵ��Gl��
�+����zcp�a4��S1r;�,�{GV�a�9W��ڰ��B��,=H�r}90��~��D�N���`6u�`��������!��<Xy�b'㷇\�NM�j�4��#y��ȬH͔�%b�0�JmN�t�.4�鞂?%�bē���OIW:�������0 �$F��-�{��w�
z�
]_I;����,�d$��bꘐd��<��,��]��
m����&t��Y����N���v@�!K�+����Z�"�`8k;z��&�V`���J�3l��ϓ:�$w�8`�-}!C�ٱ����l��V��b%��Bj������E��E���#�%��ey�}x�Vv6��r��):���K��}�.X����n|K�����I@l<��ub�Y�����'mE�	��e����oZG��`�,��fPoĽ�k�sf�Y��T��$8����D[	�X��KJ䗺�Ҍw����?�ߟH��q*25����~&��J�2���F�f6R݋�/�����3�Qkۊ|R4��g>$I�:݉O�
F���ֲ����4�}0V���:MX�_����k���`	������>������G'YG󚏃K#�j-WmqXCPd�~�@����I��wG�,V#�=�f�ʸ��u���2ӂˁb�h��ȗ�|�$�v��WDy���,^�w���?cZ�oZ�a�J�=	�MoQ5d�r?T��@��2qU�_efIu�n���7@�+�
�Nj���� �t)JY��B	��إ!�3���< ���㣾��������`ڸ(js�Z�Nb% �>�~x�}��B�U��+E}B�ږ��H���؋�xW�zr��5�����l��Ǘ�sTh��1�h�Hh��8b�	զ�q�T���j1�����;�MЇܺ��y�S*����z�w���zsp�;�'�y��2��~u�3i������/��yE9�}����0��X��!��9��b[VO���s����^`��Y��X�l�*�\[#��]m�����u.�F��4u�HR`N	3�a�	1��b�O�O^�o!6K���j�~dU����r)��ca�p��]�*N]6�"�B^<Bm������ ��wL���e��xyP�Z��w��c���M떨0|G�#ND��5��'QUs�A
�Ą����J��Y.�yi@d�Rv}g#:�\D���x�"�}�J_�j�5Ƹ#e�x	�MO�03U���5�!S�0H-��J�h�`�<_�I�o��81lN�m;G�<�W�د�"HO��`� F	��Ɲ���D���٘�1D�C͜�zg4ܚ�q�ς�(�F�l�!�M��oK�7
�����_L���C�w��Co��Z��&�L	��7��ľK�y>�C�03/9��!$��	.�s~�o�B�ѷ�nGi@�� 0���2�� )*��0Q>�r�l9�3��c7�f��ՠ���fnz����Q)?��f"�bpQ��!�Le��>�ȑ���ơL�t���9���sU��E�d�4hI7>Xݽ���w5
=.���^��C���,�Ή�Cҩཅ�`^A�즍p���2 ]��-Vt�uT)���VͦK���G�zi]���������[��܏�,�����Us�Z�=&���(��v��
ȢƄ��7�Я��F}ʰ��v8�Ŋ0Ɨ���j�'`��S�S6"@����@�����l� NW��y���3(�J
��NE��n�/���(��|����{�2$l�Ʊ�Vjy0_���k�f�0�F�<\�JQՆ�����
��yM�h��hv
�w$��*�wf���pI#Zט�X(g\�(�f^��V�t��喲���v��-β0�=�):\�mT�P�wcۊ���T�`����!�G�ou�5�_s�_�������=�!g�B�ۏq�I����x�@��ZH��'7oO�r�� B���yP���\?�"��7��8qUִ�ͫ^�b.Z�zaF�b��͐̇������,�2�)��i+���>PwK�w�����K6U?��ݨ>�0%�����F�뤙�N�ɭ��@�*�F� k�y4i�H�,��c���J��G�Z��El�V˥�|��5�T�TN�nw�WA�_'K�����+i4�-�A��T�����tx����a4D*���U��A{��V�K�H"�#��)пG����7�3\���������ga�^��h��8#�NC^��&V����������Ë��gԒ����3q��lE�N�N!z ��".�e�]�O{O�k~vE�0(7�S�Q�t�(�`�>��0O��Lb����yp�,-�Ś��Z픆� 䉢�g�}X{w�)��͝�`�g�b�Ǫ��/:R9ŕdE,����>���P
r��W���Ўɍ�o	�?k�Y��J�@G�ۂ�u=�R�,����w9���UF�{t������ Yt⁯��8m+��THfJ������&s��rqu]핂��o&����B��I�����N�����:��a��N��N;�%�B>��<�M���ţ�����1�r����|r����X�s��obM�S�K3j���z�M�[��R�,j�M�R���OX���Z��7쒯��u���e�s�(�Ms��Q�|��7#p���X�'[�<���xx�rK�D�U� !�B���uOD��Y����������2���ü9}����z[u������M���"Jԏ��A��p
�vf����L���R���N��'QѢQg�pF6V�@4��$��m���4��L�L���)'f�U�k��P��Y����k�e��rL��cߜQ�&����f
�.};OYwoUt�<�l�gT�E<��g+N��/�4�R�-/��ׅ���U#���� ���^lK�!	h�b,/3���3�bۇc
j��R�4m���b�JZ����ߑ���[�G���d���	n�AX�3�`��<�4_΢3zp>�΍��_����&�
�B�����=BVH8�u"�X�P����0�y�tY_Sx��'�}Q���:����j�
P�z�{��07�a���Q��ۤ��i����c�$�/�����I��G�6A�G���4k�����E#Α��w�=р�<�3(6w�"
V�s�1�|�*Zt�.5�O��j'c0��,$[dC/L4R��'\�L-쵉J�Mj9Y�B|S"������������
���%Э�Dp�@�\�-O^�}B���cvŀ- �u��a�o��(G��N
��O+G]_�����٪c�l�c�"���h8E��IQ|�ә�'�/�{�TQ���=į��hџG/S~�.��9i|I�\˚K%��Lo�B+�L�5�`C`�L�@���6���M!O��O;e=��pwY�� m��%]��-�Ù�S�)���W8�K�#��j=
_)W��0Uc�������%Ս����|���+�ꖚ��(OZ�-n��4bV����{�U+�˖lI
�Vjʪ��Sc��!�5�v÷ΏdR�P�X�J۶���1�B��lR�U�O% �5��� "��ɏk����jU��#6x��Ǒ�r%�]���lj�h�_�r�� ��<��O���x�GQ6���ſR!Iw�G駾�jђk�k��<����_u�,&�CŌ���P�t@p�ų��=�R�B(���f�@�Uz�ĹʗWhr���{��	���1*J�p���r8pI�u7�wen�M}���/�#&x,�[+pw��6�����0�q�kw ��b�0�-�A�����	B��k�7�{v���we��y90���3 ��ϵ6p��2Ǹ̀�Ѫd��z-��9Ś(0�.��ꌍ���oŧ�?ș��z%�Z�k��3Pd������XH�Z�ŹM2�v�����e�/;�p`����B�_2�s�V���`'����E�/�������fifvb_\Qͺ�M��{"s�ˢ]7�i�%o�![߻��/��K�U�;�n��3�RPV���^'9+�r}w���C�"���w{;�컦��b-���0�R�=%0mp�%S�n�����ͮ��+4�Z��bzG+���>(���dz@}���lA�΀�]ά����ukn_,�'Ǧ��~Y�y��h�^AeI�$�hzݮ���tYib�B9���*н|���5����]�i��h9,	H��
XI��g��g����\�ClqH��f��D�&�AvetL��3Ъ_e��æw^[xA�W	mJX��a��hM!}�_�6��J���ca�N��4�S>��E��Tg4mC��%���%r&��Ugߓ/����6�>+�bb�}0��g���3%��� 6������߰���mvk&>�}&�L� ��M~ȫ�*R_����L������i�{-R�g"��I I��Q�٥P�Xq�g����{Pt�9qa��ە�
�>�0�R��k��r� �N�C�s^F�a��%�K鎌.�����y�.�,�h�w^hr@&[�)�x`��((֤vCB�f�6�r}d�}&&h�i�)$�S�\@;H�;ղ���]�7�~�hc�	w�`�OM��E5ޔ�"Ɓ�uG����tLIrL��7�b��a|��H-�"
�y��DKN�{̝I��)#�$m�S8kU��[C`Xfiď������y�F����C��
�WG\J�V|�I�2��O>�3Q����-{ ��ig�K8�A��=������[�$b�9�D�G�4 �H�<[��?c��TK�]����L��֟��sTI�hn����9�,����+�U�|����10Y���Ws��ҨEh��S��2�����������ׄ�/#���D7S��X��E����9+���[��fJ	T�;�5�bY�}G��� u�2E.G�m�/��j�]
��M%M�,Gc��Otp{sC�X�gu؁���}Z�K��`�b��%���fd�i���,����xZ����zmإN�Җg�kr���µ�0���:I���)ĺ� p����x>�흡�U�,��]u���� ��o�!��3A�h�k�V���2�����}5��dw.���!�]�����L�?�H�Ct<&�U�D�k:�+���y��C�����Iv�co �U�>��#Y�j��o�/�p\t�=�j����j�u��L3��M�&b
U����>o���1��CR�<�yaZZ6
d��]��f��j��~-ET�aY��ă����߳n� 붒f^�n�X�g=ѷ0���Xw7u�	�ԙZ������0đ�F���^O}�AsD�k�R�]>#Z'm:�/�)��K/z3��)<�����{$���Q��/�L��O��	�t�<>�WsAb�\�w�1I�u�o:e<#���fٕ�����@���5{4���:�%��y��Z��д�j}��z2j䚉u:X��9�c�8��;>}��	Zx�%�NU>���Oս##��mRm�a�Bd�07�m�w7�i-k"��s+�?O^��Տ�0��R�F{������a�ДM���1M�A�d���$���z�%�.IE�T�:m�r���:�:�U}�w��,��@)�����d������8���z\�)$`<e,3�����pdqv��i� ���Ͻ��|�â�P��aA�>b�\[βT�j\�H;C��,.l�������dZ��M6B̶��aw�C����5��̵����(�P���,�fD�pI���-����«AL��8�.�y^�S� ��v���R��г���}�g�����V`��Ć���^#�9�T�+ot�$�d���|�>6��Р�X�_W�/O���1|��6W�z�]*:��Ϩ�����[�t����N�s�G/~�^�P_�3�d�������MG��f�.n��Ǻ	�kj,��O5�7��.8Oڧ�ڃ�	�f7&e{��a(��a:�l1:�`�ҺG�Zwd����V���r��1��ܶ�wN���1l��i����Y\d���b�)t���G��54�l��Z~�'��Hgf$�c�mN|�v,C��D���*�6�"v��!�^Se�W�fϝ��y9G͘�T��{�Z�U�jEO���'��,���1М<Tnu�ڂ�ket�v�D�)3%RM�rgc�^�%:8#������?S��A;�[�v�&�T�Iþ��`��[���éR`�U�0�G!�o��nd���l�8��Ԯ����./���_��ʅ$-sq^�x��/DZd�6U�e��	��B�/yhJ�8;�։�2B#M|$���;��&�#?s�_��gp-��&�x�������e�'B��o����Z��Hr�ce��*�T�lP�U~���nr,��ԦE'��pI�:y������cy�zr�O[K�|��kkE�@���3�x�{�Z��VR���q��8W�XBZV�Ww~��{���!�l�U,�s|���C����g@8,�*6�n���,o����#r�!���gW s��j���9��"�]�l�	�e:Ѐm�B�@g�_z�m���m��8ɑ��Z�`��$�$���!��-��
E���.��}E�vYKq��R?ƛ?��a ��_�Jݷ��B�z%B����\ߤ�^'� t�We���}�T#vvEb 4�$�D�GDY�*�vaE��B�S��̹yT  �
0]6r���&��-h4�ع��?bO��1йGu�(���dh��.��X�j J{��0"�γ��T�%�5���g�:)� �Xݧ��x��u���c�Gu�z�8V����׭�X��VY��R9���-�T��ī�"\#�",mF�'Rؠ���������*<I��s�j��e��)q���к��X9�٭?���:bLG�$l����eq�L�U�d��A��,�`3F�����
n��f̤Q�SՐ�~S#$�-�$���;dZ8��G��p�>Z(���qp���"���hF��=02�,l��:�w-�,i�K��/��>�J�F_T���U.	��V;m�l�˻~˯h0�S��{8��㇃:0�t�&�-�H�/v�&H�m������s�Jg���1ꆉV�:�O�V��l���K���3gUZ5@�M��8#:LT5+E�筳N��,�m�_�ţ�k	���.�o�4�J�<����SohS#��N'P8��s7��I�	%�{4�	�v�H��Nq��n�� �d7i3�w�,�1�a�H�C��O������$1���FwQ�x�����U<
���'}��C�bj�I��Hb������;��{ <LP[7�:
����C�HG�a�����E�������u9��ҭ�k�����(� 5+�px٫+`�3�/�3x�g�Ǳ���V�����\���	/�����n��Nd	��f�Dm����:�|�q����e�؞v�ZW�:T� z�;�q���Ē��G�!�C�̵6"�%�!���n`�����h�ƍ���W�@CL� �ƛ��n�%��u�y�AKD��c1S��a�V�-|n���v���1�|�ٿ��R�~3�@j8�BLҏ��50�����_>P�B�k��8��R4�r����3(A�	u#5�}�]�3�Rz����3F��OVT�%�T�V�>��m�ˋe���=B&wܴ��Q�ģ"6�gȑ��A�D�� 2 =z��-zDD~f�|�G���dH��B�>�h��oaD��W���p�Ev}�~�"F��
�[}� b<b�(Md�d?E�mi�p��v��0����'F#fc]��f!1�)�Ĭl��:�Q�=�9��}�D�-�qğ�B#=�%7�ۉ!h�z�#�d����)��
�sH�K�6��aD���Nl�8�H�5��lB��w����C��Lդ1�ڳi�m}���eXF9��o
L�.D�C�eR(�F�d��/=F�������%���kC(�O�|�����#���u�猭,| �^��O�2��a�;����s��2���s�ҋ���/2�Rɴ����9vF��5������`���HH���AX���_��&�A�t�l���5W�����kv����l���Fr�vo02��;�B+��et�o�~�����"lZ�y���͒��T���;��΅J��)�>7)x��s���J�U����@�F�
¾��#���&��`V|�v �_�Xg��%������]�Q�;�1Dr�Rt7��$LtD���|��#"��Q�SO�ܰ�L��"�DA�_�?y^A��u+�X&�$ǂ��'�É��Z�� 8���ĳ��C<�����S!�n闣�
�ue�ŧ��b=?��T�����\2�vC�8��v5�.�H*�����X`"���-�Y�Y�țxT-R��$  �HTAN>��+�VL�0��\aD`ؔfW�ܲ��'�������ة�u埫����Y;�*��4�ЪSt�?;֥�ܼ��`P�*IF������ם�4�%O�Ĝ�b�0)y�6C�:/$ޛV#�H���fkĕHt�,��-PU�4�G~3N�jx��G~�����:��ĺ�}ܭ��٘�ٝ��d�D �G��h��*/� }xe���|<W6.�H���<eE�d$�K&��b�����(aQ����lӁ<J���e�Ћ�ӀZ4���m��mc:WЗ��,\bT���Et�*�M��B|�ڛ�*�ܡ�+_����87E��n����GT٢�p,����;|�_5��i��'��|�N�y��ݒ��-��l�Z|��Cb����-��4H��v���������i��b%�sU��R>�«�y9f�s���\�e��!���cH���̓x6	��50�������`ͺ��Cq�e� M;��)�<��K6�X�(��Rӧ�^c����b
y_�G��hol��ʣ�]�e�{��Ʋa�������Ruhn��P8�	P ��\�X�lg
(��wO{�!\�ځ���P���2���&�U��0���^�)�k}s��u�@�P�f`-����Z�L5�2t�@�{�T�X߄t�$�Y:�<�*e�ڃ��0��!�Ƥ��P��N\YvQK�q�T1�玬7��c\����<�O�������4K-!�p�����Uˈ����}�w�A���5�cr{�}*<�Z�@�P�j�ߒ��z���Z�J-=�_����L�S0��Z��1���LQ\*,H��o���ar�h��g9w\�x��Ώ	�� �����:͵:�$�ȹ -���Z�V1�+���i��_��;+(7�າ��}��%�aQ|M���(�[����xD�~������/���:�goeH���` hJ=S�X�]�0�R�����k��3�A�C1��J�I��WHeX�L�Bn��??򺁢_ifT�`Ύb����1��5�>|m*�ه0ݼ���dkC�dn�Ӱ��
J&�Y"�YAk�E�!�獈��/a��*L?�qgt���<{�����[
�/G�<��8:�k���	2�����o���)�>���÷	��p�*\�e1y����H7-���x����G�0s�o�-!C�P,wlO�~��b�J��e��O����n�Y_q� �6�_������D^���>U��@��x��MO��}��%U;v�Bk�A	'qFg:��j��"[�t+W��rfGE�L�QZ{��������lc��.�clM�����VqA:`fR��w*����G�C�G�U��M��0�W�vŏSy�-.�<��{櫄��:y��Q�����S�B����8�}��h	Q�ָ&���Ǡk4ݯ����p�fEdz�T�޹QbL�$�W��V�-��a� �x������zpjZ1�����N�"��[LQP�OB&��Z����01�N�J��l@�ez��f��3����*��}#I���ғS�j�<��?Ea�U��F��&=^C�N���%(iN��������sL���&(�P���%}��Hm)uKC�r�*�����iJ?-��٫�:�.�ٌ�����g��0�	�s�G�7�m�mn	�cfN/<�>��?Gb����XÕ)�����޼f��1ՠr�1è�J��$r� e^*p���Y��sUf�Վ+W�ɦ�X%�qB8��ޅ�Nc���-A���E7���dV�?޶�W=��ȼF��R�h�i��䎿�h�ӥ"�>�WHO~�����$�n�6�u�L��r��sNf��h��(�k�(��_-����˞�g���Ob]�8����Xq�I�#��YNB�4��`�^7���c��4�˭� 1@ª;��|��z�S=�	����`���*q����B�+�Cj�ի�p�G�8�#Z��hRH��ގ��4�p�4��au:�f@�У����`��,��NΆ�ߣ��p�j�[���)���q߸B����V���cٰ�͂m�z^%�z�ln9L�X+҅�Q�/�I�U�f��&3�����G|���~�d����=pl���F	7P�\��P�Q_�;����d���>~��\��d���q�R��	�R2U��n�g����a���Q�މ��{�T��6ե(��Xo����������&�H'��c�Uz�m��$�}��,O�Q]ܧWpX�Go|�<4v�as�w�eEM���!�(�Կ�R~�bn����3�� �C��3�&:�s|�?P�� �bCݦ�)|to4=���3��g��}��^�|*�ܾ�]]�&ck��:�]a��켣4Ш�A�ZbJ����r�)^�x�(7e�E��[����o�L�.X�}�����i�n��h�/[��`i���h.��ĢzIw�x��Z�:�z<|#��ڴ��O���*����g>RaLfքPQ��M��
Y㤺���
�V@R6'�d��d�њ������"�㾥��
�����"#�c3S�!(�����9�5|T�x&����*w&�[�hMW �;�T�1�ļ;����������S\���w�(��f�����D���;���`�'����oՎ��KM�p>���ϒ迻zf¢a���mxùz�㧜�M	>�FRf\�BAUЈY��Z\���rR��Js&$|�`������w�V�����$�^�˄���1���ǵ�����5'`���~��Uc~"I�ы&�xU���Y�سͱ\�n�S�!�/?�
3@xI�k�&Q���+��h7
�\�Q���D�8�jg�m��d����P?93fdw�kM�ϵ�G���^�{�V��ʍF�|��ΨSEr>�m�P���	����ǇʤN�I��0P%T��a$���0����⎐}����W�@)�O}���K=��g����\�?�
o;D� ���@
�)�HC �(}ݕ�&}���Ho�1<����:�c�Bk"K���2�W�)��MR�S2�o|J*��ض�n�&�aE=�&�1\�GI��"�˫#X�����*�j��4uzup�c������5SY�Lzu��$�^�Yv��h�9zm^꿱H�4Gk��>�#2��/X��q��y�uP�G�����F��!ۚ��T�wG�ƿk��x+�~��'�E@Ap]� �5�h�VQ����=�xh�e����_� �QE.���V��E��f��-&(��9OM��>�"SeDi/CmkC\䀁?��
�7C��F�+Nt&���0�}�N�mO�v��\i�6�U����{����)(7�z|CnY��R��m���Ο'�M����"���#Z�ǁ��V�KM��B pI�鈯,�2=>ɮk�w���k�+̷3������B [<յ%�sq�K!�?�=�t�P�6��\���E���!�����|*+��v�
/]�K
� o6v�sL1!�ޔ���p�ζ���U�#���ǴW�C��j��A~.�ܥ�n-neٯ�}_�K?A�l��SB�l|Ө2����!̑��cH�A�x�ϴ=/K����Ws��蹃��?�F�r���ZM� {^�S����O��������7�Ȳ�TęRj�O�:�L�l�t��W�N]��$&c�'"�m0�a��D��[�ũ%'3�̥�8vd�nR���}��Ǽ�H�:�	���\��f��O4ͦ�'\��Mp�E��h$-Z
��¾cV�AV�d��X��ߕ��v�[bJ�g���@�����zOV�F_��墯;QA�	�+�R>�l_�I��>��p�];��jn�fP�\E��Ev�f��m\0�@�J�O�ObD:VU��1��N���5?ϑ��3�x���n�\1�f��f�+Y-^��qjݨE��<�&dl�"	~g���[�JTI-�d�~�t(����2���i�Ie8>W@��l�3g�㰊�蒖>����v<��/���ר�~�(�� �6�y\�hKt��$��s'�L���������,z��P�[�r����n��F*'BB�2^Y���Oj.��g�I"?�� �S��z�V�$��B]�����YRs�3�Y���Ÿ>jIc��%��0>������%�rm���g|���1�w'����YRo �SE �ʗ��+@��{�i ����!P�MAė�6�b���(��j,����������*$��v��iE%~B��?�H,,�4�*�ʄ�5U｜�tA:XGm���		���� ,� Z���w:�}fuȐ�*�(���SJ�=���4L���8�?�}��F-qT�9Ε�Ҭ���n�MGG�*E�~R��굾v�'�iF�+����F}���a/��"s��i�-ْA�ry����鋭η�|R��lW}V��Q]��鎸&Ő��o�8>��k�o#_�+���$�,!����$>\����[/-�r��&���y�:����x8RI�l���4pN���}A
��޹��;1�]�[�ތ�:��-�V(�p����Tը��j߮,��̫��c�Ξ ���n��h�F��a*�F���ls��w�$B�M��{./��Yi��5�`�D�~\�p#x�7Sk.ǩ�ĕFr�����������T�਍���s9�f���]�y�h��!g�I�H��s����Lx��y�(L$)S:uBzU`�@h�"��7���y�ڬ�)F��3��^}RdpVy|58��T��;�rc$����l+v��τYA�;�5�u��rҀƩ��&����;Q���nk�Ǒ=Ձ��P۞o��9����]l����\F����4�s��i���{�R�
b%��9b!�g�:�QAI�
��f�꒛��J�X�i�W���G=�XX�Y�b٩��n�T�߹�b9�ӓ�0wIǂm��#Ʀ�e��3h��&�׹.?Oб~���g�͟fa�gɴҳN��ѵ�t�Ϋ�0JA�ǌ���L�6.�H;5d8o9갷��s� �|�eF�%@f�3���O�p
�����ܙ;Y}�t�2��}9{
k!���O#%ͣU�A�Z�~��Y#�1��9���+)��" �y���*�d��h��"�Ɩ�Һ��_�Ȋ�����g}eg�z�K���Ŧ5i?a��4+��&�Ĺ�=��v2�h��?ٲVe�&�ⷼN�H�ЏX0���-߻L<�rʋ�W�N(��kӡ0�xΑ��aU���/�&w8p�~��7��:֪DzК(q�jT-���7�2M��xb�ա�e�sYz�m��̈�d�RX��ѳD4�4��o�bnwiH8"���XƗ�����S��+�GcDy�LA��� �־�N)Wm�"s��'Z�T��1��)�=i���|:�(#�%d���h#T���mt>�8��-.~愤<�r�\�*��Qe����σ�&���w���H�d1��������r����j`NIR�:u&1Q��M��cDgv>o�%q-(ţ׏[|A�^HP�E�E୕���J>���P��Ǚ8�x+���
a~�lH�4�Y$�����Xȥ�z� �	�\;U���١+V�gyQ��)86�{��w����\��,�;�ޝ����xP^�3�W���
�D����J��J���M�(��U��*QS����A�e8���_��9��訞w�a�-���x���raa+�Cw�K&G4-��mN��a��r���cH�
��;V�@:)uی/�MI<�䈀R��z;dSa�ʕl��$���H@B����w~
YQ�7��O$���xU�OA���b7�C�uՒ q�Esrҽ�V5�V�:�;l�'�F�Ӱ{�F��>y2��}�e����	�R�z��Ě1%�΀}P;XAW��C��[U"1�}�K�6R������w�6��H�ӥ����q�b��o��#��X��r:(^.pt���R��A��$5c�d��_�j%J�)Q.��J��)��/X���f`��پ����7V*.'e$<��,$�XKJ��c�a�v)<邾����`��b�GY;���i���
���;[4{�ף����:�$�����t:�̈́�+(3�zU���E��@9��O�E\r��R��S�ܧ+�~ �N���V�X��L(��Q��w��t�0�ˉSE����p�:��`��{�m~]���{C�U*Z���.�7�^: l�R9U�~��!C`Zu#�'����Ĝ�0���� �����E���c|`�z<I���@k}W�[���U�T�N�<�af!��SNm�4�t����F�!��`軞V�y�Z,b"0����6R����დ���V�1ר���%��9ֲμ�l�spv�RfC d�%r5x�J�7؝��/�c>~ ���������/Υ|�Q��m֯��t���Q�<�>NM��i�{���Q��������x��] Kڟ�����~���${_�45ND�z�L�o�ط@���5ko�g;sׅ8�|�E�4�����|L��H@;Dl)0i�p�-��MY�=Jo*�^�_xҮ��c���
���R|��Z�/�(my�r_>I�B�74e��/y
7"� u8�i�U���I�����Ofs4_�3"��7�w]�׮Xs��f�,|/o��̺0�����U0��L��?^��O&؇�g��̸\X�SYDG��RS��Μ���Bm�ݭOuF^蠎�1hZy��TO�����U)ʘ��-8��2(��B�-�+���A�6�SR):W<[#G$"0A��j���~㯩!�q�������8~G�Gj��)>'��A@��!��乼#?)�ɧǝ`���>��S8.��{��@/	�c��
l�aA��A$H��J+��z������e�\�8�]w2|#��¤�-$	��JɲGy�<cl�ب��b�^����R!�#���W���!��g��O%.�	D��e��d_j[}g-�����<7j[6p��ʊ-hךX�����܉���s�[�G�rh���Q�`ak������y�g�W_�b�Y"�ڡ'����>�;���a۬�����ʉܚ��?���A��1�f>2�tR�q�&��b�F,q�%��0Eh3�n��WlP�֗e&f���8��Q�?�t)B�}"	/�,�b'��G���W�g���$�h���ݮc1o\�"T�[��I/�>��|b%6k�Q��	Ra��V��:��b��ty�p���[���i	2�ޝU��p9	\���	,�ו������9d}�
��:�c���z�r5rܮ]D���kz���ZE�P@�؆����Q�4i� ����s8n��sq�Nv�R�Y��|0��@	��_Ώ4/4Qf��؄�S�R΂�I\i/�9yF��;XW6������	�\x5�߈~�y	R:-/����;x��]��:��kE�yk�����������T��)}�rݜ�of��΃�%: ����9�@�N��<�M!�!ٻ����-e��~��ɑw2�i$�a�h:���Xvfgݱ�
�Z���\kX,��;���_������	�pj c�N�(gd��	#b@?�(1���|ا��v�[�ӷN}���}���$��o�
�^���\��/���1�/������j�n�}sq?�S\��x=�Z8�+穓�����@Gd[qD��ӯ�&�\�{1y�@@�Pup���č��������
��O 5���o�c��� Ԭ��m�I� w�(0�yˁ�����։�5�z0�$%D��$���Yc�b �e���M�};�%ܭ�W�A�6?�T�_ �a�k�D��y�o |J�r����e����1���%����W{Wh1�'0%�c����o��NJ�:�X&�^[�2��(4â��E5�/)j6�D.�$�am�dS.`@w�O�0���6
�j��|�@?:E�V;�(��L��h�zD�g3B�N.�e���B�:DiQ��D�3��+M;B��Ж�1��Q� %u���B��'�¹�o�%�*�l����8���y�AM͛[F���K�auS�z�xWL�����Ln�c?�U=���Di\����>��Dׄ���W��\F�d8I/� ME5(�`m�M���7�FU,�����f��X��f�+���o�rs7���p�.f�-Nn��y�&!��N �Q��߻�Ť�rP2��^mD���X:_�c⋃(I�M�X9�2SKjS17�9�&0�gq�;y09�NXKs�/؃�[T+�ɾ�%�Rla�aq)��r��E�m{����1`���g*��/#PT�zB�Q�v������6,�U��m)/ W�^���\17�[WAKv`h�}�-Ƹ*tT���y�[n��n��˹�;XS"�q�(�u"��r~v��Ģ���Nw���k�u6I4KT;8�f��&`���yP��f��)E�����T����2_5�>���3�{n��ex�N�k���sx\Z���%{���o8��N���u+y� ����>��h�H�S!Yǭv읻POn^����\$h�[��j=��q��$�����x���b�>u^�~Ќ��������Df�ק��l�[��lK;�)��M���4s�q+_19�޳'_ק��w`��mZ�\HW���P���W���f�z�)��"�|����J�F\d�H�"N��nI�(�>XI�PQ����س��7u�{�������g�v ��{]
�x�`q��~�����R#E/�i)��B�M�����tjZ׀Y����r��S;����>-+�'�F�����l7��E���(���{P��7�<�N�%���(�mB�N ���C�(�+�便iS5-I+�3K�U�G�a��[� �X��YOz�?=�#<[D�#E��;��-����O0��$�ݙ}˗��`AR����m^E|<>�� ���� [�JNs8b�Y��Q?��,��w��"ec�O�0I�gh~v簂(��`�*�4�'gh]3F�f�����
�)A��=��}JTGh]�� R���4Ά�]��5TJp����0�5��;�Va�ك69Ex~pM9nͻ�����1�N۟��	-#x�|��`�[k���� ���I�i��c^/jH��%�&�z�'�����`�d�}��v�����b0Q�Ҫ!l�ޫDx�5W��h?������X)���T1w�)*��T�7���;g�a���4��`Gt���ژ2���x|ӷ�i#��Q���8D�g�����
�O���i�&fNo�_�hM�����#1��xE��}v��`��@��j����
�<�_�:�f�'��-.?p${��x!�SG	���������9��=6?�&@+�?v&��_[��*���%�^�	���	gFBK&�U4��ۨ-k�?��Oa�Na�Bm��W�F��ه��9&*b}�砱�]jMa�u��:���,i^�#U�� A�?�o��p{ňA���B?�69��Z�H<D2����T�k��ꝼ���׹�}�%l$
\��K� 蚻k8�xh�	D�+��Dc�)$⊩�2�; ��84d����sCs:�P7Zp�[3��)�c��P�h~���6�G��8�F�j���������~�Ը�TZ!�l�Z�'�E�ZL�=m��U��k���*r8jhG�<!L��L�t�H�*�'�'��	BKo�2��Zh2��E�Tȡv:��K�����=d�P�qkMՇG��֫\?6��@���,���¶�}�1$[<O�(c>�4$o0�CL���脾t�n��n�0D��> �v9[�#�O庘��%w�1�����gGU6�f`�'�6��_�h��&O�js����B=M��1yh�j���5f�������c�f��l����A'0)��׹1�G�j*��o8@ǹ�t$�7�-[�OΫ�<���ܗ�L:�H���xġ�-`~��z����S���2��-	�Or|��d�r�I�q�<����u��ܑ�v�+�[}���Ny�������-Vn��U8._b�`n�6Vi�����������o={�yet1�;�y�Z�yЦ:f������9�i�;'�����Y2�ӷ�Y&C���dk��%{f��o�5�n��\���I��7��+V��E�.�z�	��W�#���T�.h�l�iE�X�2����.��]��XϪ��k�IډX��Y��/���8����H�g�k�X�v��3�C)�7���g���#@f*Gi��ɴ\���s�zI�Z��-�8���f�[d�rt��E��D�20l �QL �5mpR��!���`��B	z��Ӊ��j_s�Y�X�b{m/�v���4�G+A�,a�H�BE��_�<�9xv�;���0-#�ı @u���U�
q3��2�h�^47�T���:�糣]�5��$9��(��Y�2��K�U�,�tmd�숪���߮��n�gd=�.��(>×�&W���0:\�.�>�du���K�dp��BCP�u!'M�n� �H��Z��]EFtWժ��|���Yr�R��2Vxh;��"9_m��(XjL��%�>��/�KQ��M�:?�H�s����4��)�� o��bp��/Tk�av��%7ݿ���6�zm��"\���L*+'�v긷�C[*C�������Ŭ�J�r�@S��lX��~go��|
L��*����Fn%��[{���b��G�
�	�[�.P��Z��$@VL�JkD�!~�:�nŕͳ5�4��D�!k��[�/�;�ݦ�Ϋ0��Y���
�
W��l&7i�q^r���⢷��9������v��`�H� �w1�j��.�6(����(�zd�G]{*-9�CS��F5mC"��n��������S������(*�_�*���֘Z6vzf��5��B���ǂ%^6/뺒��%�.�\��ķB��>�m��J���g�x�2�3��ρ�d������B��C�!�yR3��g���9eVnz��r\�!
���:\��[�0�d�!��\|ٿ䜳讇/H>v�)>z��AT���H��~@7t��S��J]����zF��c"���}�K����p�������h�wI�[/u�}�0��q��\0bx�bÚ��	P��( ��c���B�p";y���lE�	�%�J���Y�������;��	fO��=n���,�.=%��0u6�	����]F3x�4EQ�z��T�E.�-�f5Pt'���X���Ц�vE���u����XJ���a�i��Oa�Ӌ! ��$'�E\�]��,������S�Gwscl��5�8���/$��E��G��w�K�p�}��T��ۻGV�����(n-�^e^��A�r֬h\%�f�Y���)�dt��o�9���-rU�z�u��Z��c��hy�s���-���7���UB�(������]�i�j�J��q:�G4g8�֮�g�S��8�Y�&��i�����DV!-�h���u���.�j��,���+Q|Nǭו���vmO�f��[�-/ �?"iu�5�r)�z�>�;�0�K���zW�U���J���J����v	N�'~�j�M������&��$���Q�ԓ �%�)�X8@�y�k�^:�B��+zw�V�v�֞m�țQ�z9�c��S�R�:ţKL\ʰ�@��a-�+��j[WQ�D�2`�R`��̑�L�����~ �F�_M��HY�����AA�7�Rʒ��)K��4�s3Ƣ�j�:��C��p�/�m9_��&��I��د������uN_�<XS�V�sC'th�w:��({�$8C�l������=t�ֶs����?��Q��rxYL*�A��<�}s�d���,�G�v��5�������[�y^P�j^�� �B��\
^���?�<��{�$o��Kb�r��fLF],v|���o��E�������p�K Z+�!&l�CZܤ�q[ԥ�ጙ�Z�m��|]�t��|����x"�R�S>�"�Y�Ayw%+�5���do_¾�����ꫮ�������ˇF69�W�����H��޴W1geB��_�AX�&X��wD�	CQ�MP2kl��Ӫ����hI������ujm[14���k9���̖yd�AV�
�����{xuM��q� ����"��
Z}��03��D�k|�r���*�n�^A�������a#W�n��ɡu@�ظ��C�C?\�"`��˼_���#��i�
4Tz�N;�o1�12�[	ԩ|7�����F�
{�I��V،���1ȗ*V
������-��3b֬�;�[ ��> �*7�K�.��P@��7�ΐw|H(�|��(2c�Y{�=�M��e��4���Q��"��²�08U�I��z�s�*����X)�0��3��=JvCY��Y??zBT5�5�v�{��ٟ]!t\�7�DJA~�W��l���� \f�E�����r"P�r� �g��ʻ2/ѧCs�G�-,�r�J
*���Q�,v>�F��������gB��GԲv�i4���� ��Y<�&��by��)���8<^��<�5�TJ���BS_+���M�oR��T9���m���?ZG��A��9����`�-��An<V�3Du�	��.da�.��ɖE�=����/��Kg�4A�&ͻD��?�W˔HpT������V��b���$��Z!3��$;6��&�]ѱ�{��Z'���4�m\�E��w��Ĭ#pEK���qB��d����bx �,������PB��M+��/]������R��GA�c>���L4v�z����'��X���1.j���*È�g�5y ���8ji!�dZ��m zXUӧ��#��;���bX�5��
��z�m��!��`>�v�<0����/�������W^��>��,�K��+��������Ϗ���SX,R�O����.D_T�r�Y&+���ʝQ�1	i=���I�R����1}$%��x�?���3E���������Ek���l׺���Z��Se�Y�ę�xG�R�2FԳ��\��Q�·S�O(�x��񍀥
m{�e��-}���	!\G��e2��!o�?QZzYHA�a��#b)�j�I��u�I�qw���Y'a���i���k����G��w��C�Q�aM����!���\�˸��0��5��uO"\?���R3A�L�"��!s�+$l�r�A�̼�&����m���X;�`>v~�7���Ss��J�R��]�a��2� ��X��R�X`��F�xR��1W�m������!�� Q�h��Ɨ蓺�b��;�Xw-8�,k^��"���� �G�u#�*WiT:{�)�56'?�jUL#���;4���r���}���_�.JTɯ=�Bz\��:���Jo'|�@�P�>���KB��b�Qu#,n=�=����Ùi�('v��u�#��P)���?��.B%�H�S�E�Y�g�����9��艰Y0`�靸 �4�l�;��K�E�{����f�6t�� �ܸ^k���^�A������ޛ��"�_�3I��1����?q ���|~w�Ǿ��gn�΍���Ţ{�γ�c������\�|1�t-���=40t����j���H����O��D3Oj�ȏ�H$�x�1��]�s�����O���ϫJ��5�~�����!��%����ܵ�y��NF.]D�2�20�6���F�鱭<N�]rpךt�:�,��4�⊼�kϺ)�K���ػ�טV_��W���U`/�"��V�0���Fz�a���q�tc�w%hx4��8�,f���:���8$��N�J�j� $��MNA~���`����j�p�;ADHM�(U�d%�.�#&���TI^w
7(KN�:�¨Ln2.�-"��p��Q��2y��$����*6X��Ԁ�C�H�b'_[�W����k:�p�'�8׻~��H{������C��d�Y��� %ƽ>Oz�e܅-�:c|?�rM�3/��'��MU*�N'�[ˤ2Al��.�X2�3�M��F
�/����v�io��Q� �Y��d��-��X�gR'4&�-
�l�o.��.�"sDN�K/B+9�Sl.����������f2����>\4 Q7�8���ҵ0c���R���J.;�MP�Kn0(۵M*/��a�}j���o'���c8[�@�f̝�U�Ǆ�e<��*�%��,lg�h}v���q�]���c�u�^�([��Q��1��CL��B��A33�5<>������dP�˻7А���7H,^Z��JT�+�P��e��N�S�r�w?��8����G�w(C�[Yy�-x�-��st��|�ќӵ^g�7��z� �1��F.�bW�q0s��ѫƯ�.ʡh��A���BT�*���WA��Ia�(�ؗ��&X-�L���7�<�! @؇q�[�r���#��Du�N�Ž�	8?砯H�2pk�Z�A��Y��C��/��Yi��G�/�n�S]+��M� �r�h��d�$�2ٝ�`=v*j/�n���Q�P&�I���0�@d(�%�Ö/z��b��^�	���2�e�ɜ�ĕ���q��o6P�0g3�U^��%��*DV+V�_��Z���??jTiۆ�����t�Yо<��1�7�8^�/,�".XF潸��80#J&m����{:Ɋ�$ud9���E��Z��U��'�8:jK���� "8F	��f=?�2�]�ǭ�p�S�c&$E�7%G#T|��Ԕ�
����ۇ�f��:����;�cg�»��h{F��[��K�
5���bv'�wA��a[g�_���Č��#�v8�eѥ�*�GkB��Wߛ�cJ"Ti{�y�V3R�F\]���S�Ћs|�3�̓�$@�֊ǜkfR�2����U�e����-)0:��m)�}�&��C�(&�6md��\'�x�%=#����Pp��,Ő�eW����lXz��H�>cB�\?;'d, ��O��Ok��=5��עw�,3泄7=C�o~m�HP�nz���MDtGR��^e��
ݞ��Id�!�i1X����_\e�k�)��ݬ	�}�	V��<�g�?	����O�Il�A�`��	cx����;b�r���"���*\��u�Ti�߃���� "�� vՠR?��#��f���:D���UO�S�y�Mۃ���QQ��dwx.Œ��Z�0�#Dp�����L��30;!4��D}�U>�0�.�T��i�Ž�b�����f�P��M�;5��Oc�ݞ��O�:F1$ݚ�I��hC��I���1�J�lpbhR��	���O�eW��㐔-��&AE����}�Y�	ɳ��)�q�SG�����K�of�O�h#�3a��b��Y؆[�4$�8�u����z�($I�/�E��ɕͿ��H�_�4n�NI�:T���B
 �1Q�P�b�mxs(��Hg��8��CϹG��soӘJz�����t�i�<��f��c(���%��]D��dV�-�0�*53� hw�z��^���e��.ŚeLfS�Wc^7@���SK�aGs���&S�����yW�䏽g����w��I�ݢ�e��IP�V���M�v�-~�iF
�_��w��|i�ś(qQ'�x9���:�vAM�O5���<B᳁kI
¦�H ަnJK� �����lM���-'�̟|6��q6B�wj� x�夻��:��jf�0LǙ=�R]�Ǉ�=�����w������2jʜ��>���{j�8��C��ej�j��L5���g�����q�J!e�r��D�,X+������'G[75���4��ğjϙr1V��s����̣�nJЖ��f��0�r�^�0�U۹#�WD��qz��цԴ�� %��P����,����7�qt���Kk"/�C5���5�ss��2½�Y>U+ ڎ�-�4Z��y���?����AڊSCLA̭�E���P����G�����9
�?�H�$�Ͳ��`ї�~s�c���E���?M7�)ț� ��8�xR�'���_���,|��B�=�*p����4�B�j�vm��ʚw������*ȍ����T�7����#�*�b��Գ�q�F/���cܖ���n֎� �-�¢Ȑ/sU�U��H��^����>�P5o�*���TG�VL3fl�B:��:��)p���`��:��<��B�5���&^���\7L�}hQY+� ߺ$}�H�X��!� I��a�j��M��x�b	���b/�ۃ}�f�9�s�5lT!^�?����E��tJ|�I8��KB��D�fČz�f�0�/�PI��� ҋ����U���*���ߡ#���
^"Cr����;i�(���8[�0��{�	�ob9���0�[k�#����`{K���րl�� u�!h���r�h���hbB��Ln'��؋x-oHm�� �6l=i�H�j��%�y������u�ϣE��S�b����"xj�jlU��)Ly����S��a���7�v���|V�{n�hz�r�ʃN�}|r��&�
싌�iޖЏ#�Z TX��||N��64�Z����ۃ.�4�z���Z���NZ��p�.���U[�S��N���=G�g�K�$�v�S��k�xl�J����)zr��2�T�Ie��t�@t�0����1�+�4z�*^�<B#�5NW�~��ܿ)�BI�Z�}A�T-���M�I�'sh�L}�Q�hb�uZa�������/LUtU��m����B��T�ɧb�o�OHಯk���������0Zo�^KڛY�!A.-;QTU)l�1>�~z�/'�p��o+k'�8�	8�ﺁ��og{��U��c�T�_к�"�~��!dA�f{O����h��ڗ���
�"@� T�U:��&Rb�ֻ�j��� �n'T�r��ԍ�Z/��S�`K =��kP�\{W�\�n�<��źv7�\�Q�UG��"�>nhQ����"��ϥ�+��LhrE\�����ka�t��g���E����]Yp����d��8"����Ӟ�d]����h���9#�����?L����?<NF��<�嘢+ٰ�h��N��n&i����	����ȮD,�S_���#�,��iƩO����67&eלܭ�6(���0���뱥�򍷾F�I�rWj���P�jY?���c!OcD��a�'�sd#reF��H�����w0�јk�:Zh���N�GI��Q[�0&��:!�ͣ�8Eu��P�N�7�s3����|B;f�#,߉�̬�|��P�=�4���Q����2eM�lPU��o��^&��OI���D���1�@]�h��5�ԡk�㱲S�����B5��D�/p�5�4)�Ы��~j��݁�vS�X�e�d�E�E�Vs,�������T��Ɇ�F�g���9R=Oj�k߁��e �%I�^*_	 �c��W�b��:�ߴ�h�	���������0R��Ϗ��J�ϕ՟���)��yzX��?g@��ױ�����Y�=�Ta֐je�V�5�֑M���+��CZ�"�e�����Q�A �GW�_0���5L����x�,`�����?�H�X��7h,h�������Kڭ)H�x^�������F�g�(�E,T�k'3���W�<P�)�K �1���%/�!�o���� �_���<����܅�a�֝��!\��q�D"C7yZ��n-�r<��]oۀ�n��Ʉ#�WD��h�B[	j:�:8�����y+dVF可ԗ�8!"ھH�\�T�m�[,�w����+�W�sr��DuWy����>8���v>Z���Q,o��.�aG2�d�T	�$��m�T#�����­�
x��	�d�#��E����$`5(����OG�%2�3�;������ĥ �4ܦ޵�?��U�M����� ��?�"�`N�5�JV�&܃�����&9���*��o���jM ��m�qy��h֖�'�6�e8.���p)7��U��v��>����<�:��� �j�YT��U�mK!	jVc�0Ì�5�;�6HQU�����K�!�e�Q��5��P_���9��ݥI�H$�"b0�n�������X{��ɂ��� O���K;�T�t�SI|��a��v�2��x�V�p�����x�n�r��wE�N���1�Q�\/?. J-E�xn���x�{�O ��\��ƴgm�Z���Ɇ*��1�����M`�7�z']d*~͈}���q���^v{y�e&eؽ��pF#,@$9�ÿ��ls��.�!d6 �4�6.�l��1b-�f٣A 9�-�M#�dvdP+t`2N�r)�R�48z�2��im�{-�jg��N.ʺ���4F��1�n"2����_�XOt�&�d֧��:�����j��`�㆘c�͞`	��?"v�'I��IG��i+)<�O�?���<8�6���
o E�"��/��НI%0����$/�Ffp���U�`�����&{�.��E+& 򖍢#U������M$Y|C
c b}�n�4�o�`� X&�#��ˍ��ʴh'�otc��p\�6��#;8Q�uA�l��px������|O��
+�r;�+�g.��P�)v
i�NTs5#�E��j��d�K�L�.HV�ҋXoO�Z���tř;K��\���\k����^)�}�-�z�-��0p��2�E7Z�y��_�0lN��~��$��e��Y#{C�"˻��ge�f��d�V�����يw���`���C�M�8�oo�I������Eg����ǆw�K1�l`cO�<�|Hݓ�+��]Iէ�����2���V�҇,�u=W�ф��e�<�������-�`�F��{�	� �s7�&&)�lh��'�]�%�7 q������d5m �� .]�ђ�ڳ��
h�g��U3��N�~K�"]\V�ٗ*�9)��^k[����F�[�]�(�����J����Lu��z��!U#	w�4̣���p�d��~zM��֖���Ӵ}�c���7����G�<��/#��6-��.ր���;d�h��-ʯ'���]G���\�־�i�e�������6�C�rg���f�E��%}Ab%C�)T�Fg���=,uL��2U7�sC���%!��~�K��o�����,��r��6���
f��Kg�|D�\�q>3z�{R��̃�d.]�|����`�yP)9�Iq��2����e�M����If;קe��ZJ�6pe�QD]��p-�۔��B̦G�uZ��XzoFhd$�'�W��^K�����8/+A��=�n��c=#;,��$�\^E��XxF������2�f¶���&��r� ݡ��(<4C�+��'��ޓٴ�"|��ŷR����Wa!����8u$}�\F��jW��HS����)l�-ݠA�	R�>�o�h8(�lvofNg�D(�d@�~�6��N%[�M��k�x�ﰣ�t���+LT��{�f�Z�o��\�V�b��ZX$ �YT,,OU_)P��5���t��j��><
bb���0��;�ϡx���cZT	;1���;R9�i}�i�v�n>��ɽ2�����w@0�+6�{�r�z?�x*T���_��S�F�K��b��`�Bwa��H���	j���
 ��Z'5�v,��)`�u~��,������H�R��2J�"Cu�SD �AԸ+��!{�����0ʭ���sF�����˳ ?�[�Z�V��o{n����[��� e�<Zl!�������/��̹��~:@�>�R���B`�Z���9:�=�C������ß�>UGz{�N� �!����V�ol��6z#!� �szS��'�-^�e�>�S�V����\������6Id�g��"�Q�k	����f#"ٙ@�����o�R>�]v�Yy9U�����q�G+�iKN��ot���&���h*`}��gࠡ��K$ϒ��Oـ�8Z��ܹ}�:ֽ�)����Qw����iڋ����t�{:�`����<<>X1c��ֹl")�8����҈t��D��t��29�%��M��}�,���˰�����u��U:a��Ƿ�$$.�<�<��(�!��
/���k���v�Qu!2Q���/c)Vx$u�6��S>
I.�҄YΰF��/[ׁ���i�ta�˙�� f2�+I ��ap�^u�C*�\�c�FD��ި+��/BD��\���3����s���I��c8�L�[����P�E(j��~􌻳�\v9eb��ˎ���'��,����k�IplF����P3��>I(���� 	�p��tgP�:H�ǆg�Ȟ�y�:Q0��C��ƣ�L���v��V��9�ן�ZǞڠg������bT�������$��7m4����x�I�T�6�4�W�,�p��72�i2Y�;��<x�[��(P$:.=��1ʄ갍�"l}C>�nc5~^����btG�>�w\�n�1���[~�T��wT90����F�P"	��e$�?��EX @}ӗ��]�ӎ"f���x�Q]��9.���o�)�B�פ�#��RKz<�-�����dJ]�]��r����y^~qC���E�13k�6Wߜ|�]=5y=��l�����[)7�`Pc�̤��~9�k��j!����or���ը8��) d��^�5���� �����<]�$�<S���`��Չkٺ��Su�4��ڐ7pd>��(m�F���=���+����T�.6��Ֆ�dg�Y�*n{��-�>S��l��̐s�[W����o\��f�Z���rR]����(�����k$�J�2P(��d���������:��}S���ɸ9�Ĥը�r��s���x~Ft�Pbo�"��>Y6X�V�}cJ#�����F�k�|�0'�Wh%���
bT*�PC���V��L<�[֢~.v	C z�j�psSI��+{7�o��|�W�̼��a�,���5��?�w�D	�R�w!��������G���B�'J6�Bv7s��E�|u�+�1*�A�.�WXg(�>��vV{�|Âؖuy�{DV��� /��b�T>���ߪ���Q�Ƌ�{�MәWĿ@�7+�����p� %C�ǲT��R�T�;�yY���Ǫ��fJ[u!�r�d���zg��� Dv`U��['�wې��ĐB��嗟7�e��SP蟋�v�.�J�e�f%0g�?;"��v]�`�3I��ovC�{�U�˕W��w�(+��O���<�(�7����R�,!?���NBeA�6�P�
�)��P�1�Sd2�*{��6�Y`���Uё����˚>>�c#��m��Y��Z�{���6x�z`B��)��j%�� �sl4ػLD��D���;?1�C$�K��Ex���J����ѡCY]h�R���;b��a�k�� w��Gg����JMj�-��aK%:F��BD,�<2���|]:ǧs�1rGT�@�Y��6u����"q�n(���9VT[����;���0<BAN���D3̃���B�/^^��Gt�Gᦏ�6b0d]Mm��t�:��q���t-�V�J���&'і�H��C&4��B�����$����SB.���ߠ������k���1-<!�{L�R�#�g'z���$����|�TB�,�O_�!@k�?,�Qa�ٙ����f������!�ԍF�j�f{�& o�ig�D�̵�w=���c]� A�V=$�[�	*EW5�u�ffq��<��֩�x=�ӎH�y��ņ�Y&n��{���4Y$V��_��Կ����=#���z>�4�]>������KuV��6[�[|c�A�"���o�>�(�i��G��t����p����פ�����/߉2���e�����'{vC�al�DoA�\�5H=Bv�W
��ߋ��w1��,(�!��JQ��2R(�5֟��"n�{&?�)@���K%����f`�@�jfC�ܔ��?�w��D?������_tc[�7򵑰�~7�/�	�	���:C�}C�Q�j��-ͱ��E��*
ש���0_:���#��
���_���v��n&��������Z�R�h�Q�*#k�Îş�n߼�=�,R�ԑ9���e�����DAX���ŪK�p��,f���w1	j�E���7�I�e".�V/���UAE9�e�2�������"� �L�c���F #�n/��Ky�6x�mKW�=}�|F��j��v����Ib��'C=`������Z�D���d��]*��a��ኙ��Wq���U2�Oe���|؛�.}��/�&���_�v-Ƌ�Oa�L����ns��I��fG�.�B-�Ƽ���ס��^]�	y����T
0ݏ脇��	E��2dW��j�E�m�j�b��2f�J�!K�.�$�{�w�ߊ����Kw9W�@Zt$���.OQ�$�ëU)x���`2���OQ�1Q��R>���=�d&)_J/�R��d����2l8-��M���k�w���R�0z83H���+��L�Unp�IX��e�D��Ј(#�#'@�F�2y#Πs�s�Y����r��.����#ξ@�y���OC.�.!�5w�m�[�r�;ں|v��}��O�>�)�T��a��=�u��d��j^K:魦�X-�����C�<�b6B\���Z�6��t��QZ���E$�/ч6��;n&f�w�x�T�,���VS@ወ�J�vN��V�`����͏����!�V�Ā|#��l0� .q�~�%��x��J�h�����u�רb�ص\�|�p(_!,���f5��ܰ��<\�\U>~����
�>Vo��5D���!���}���AVH$�縫/�y&�}�qh.4ʏ0�[쾈nY����'�<�v�:S������W�v4��|�(�X�߱A��bX�;a-��*�lg��'s���lK�B<ٝV����T������6-�I;�>IhV���3����~.픶	#���P$�?���2���z��c�k9�ķ�An���=ʪ�'�%���ř]^vՒ,Y�B�5[Ք�w1����5Wm�Թ��`����\+��㗅�7��́a��޴C�3a�y�`��� A42v.����p�X\R��Я��`�$�u�#�~l�Ch����M�իߕ�`�(_Z�ڱ�
�-������m�ٴ&�͞m���eC��rH8�݁Ƅ�#�'XE�<kI��"� ������Z	�����kPy�(x)`^.��"/�(���q������]Ķßd_�B�S�?p�q��Eس:6N>�N>�W���n�`���~��]�K�D�j&?g��p gd��޻:A��e���ݠ4�z��!����%�.�{+�d�7V�h��Pr�Q�ұ|����g��k�v�p�$��O�iM��&�ʷ��5��4,ã�����h�=����SO��X��Q�)u츰,4vǵBU.����&_]+�&>�A7�?�E�
�$���"����(�Qn(�g��d}��[_EXEF����������/�!E�/�W�u�Bp�]�zب�O� �B�;�T-�5+��'�v�D/�#��U��<����3�-��D����!f<���i�9�~[ǚ���.���.�jڜs���S@,9���SǮ:�E]������4y�i�����t�e��i����[a.#�ܭ�v{ѯh�_^��H l�	�/��B�h��'CC�WX����u���d�Q��}I� �7�10���?�06��˃M����Xޥ"�ѓ��a��8�z�dy���)�@���ˋ7T��+�.*�V��h��V7���*�ѓˇU} ���73�t�H)9]�l٘s�gBY}7M��Ǯ�F&;ԑLA9{a������2�V������2\�Ԁ�~�q�ժ�T�~���%���3?���ߜ�3&�R5Պ������{�#V
� ��I'��< k~ߥ؁E����aV�2.}�5Y�I��C�v+)6~ž&�-a�� k9��a!1��� 4%�Q��}���c/LF�i��NB��A����7�%Y��oF�㩃d��pgܸ�E��`����3l�Ub%V��� �M��9(���������p��d��<3��x����ء��1�X�N ��\c�I7�qg^m��p�n��Op�Ԡ+�� �[VϬ6r+�Ĥ��[!��n�r�3Z����U���_j����<:T�7���&�6M�9i��.���6=��:;�y���9���Y�"�RG�]n��k�9
���_�8�w�Y�U��p633Xqٶ:Y+ܠ_^"�[N9�օ_�'1g-��j"D����tV�~���z�9��q���<e��v�KL[��=8�v�1���)���z#�4C }��ȣ�|�?�d^VQ�O��(��=�4F�A�=���s'@�J��8aȸ	�I�����Z��~�������~�sUs=|g�d�|��>ހew�h��^;�7(U@�����'C�'�*�rה�����h�D��/}�2�}�Y����<O�*N5G��E���;}M��7���>e}�r<NJ��*6�%0�o��a1c�, U3bQ�uz�b�}c�Kw�<�����z��i}��>x�ʎ�؆�u�������Fsߣ+|�,��t�בA�+bQ�9��p�:���7pW&$L]S�a�L�aR�,%���������C�����AJ�;cƹQ�'lq�oh;�@4D2U�ɗ6��`y	WD0��!��~S�fE������QH�j��x)�ħ ���aY�3���YT1~1R~S���>�|����GaT�j��)U,OSt�������ט�{�qs�<��{�ޫ+uP�uI�Rt�~`o�����X�'�BeQR�N2���� �� �2�8\�����7��)�l��!ܴ�UŇ���x�ه���"ّ���K:ۧ�m���R�(-��;��� ��B�a��Â��p/Vc��!�����ʬN�H#L�b�m������`r�2���� eޅ���3(@�R���%]�SWn����ִ>X:�.�Agͷ�rh��X��W|��{y>�&��dP�ٻ%q��
;1���i�������Q �滑d�,���1aʥŋK�Y--�u��euv3}~�.	.-j_�e�2�������?�u��F=}X���;�L��B�����@t�-k=:��Fh��_�l\�A�蛩��D�ܥ�x�JH��/�t�&
�������<`\��=%C�P{�е���e������x����E�b�dא�1���S �A�*�����rb@�S�Ì��XN�Cam'
�"-Ay��A��:Yi�F}E[5>ȯA�����]H�1v�p�ca�t-�|��`�^{;ZV&�>��E�'��:8��C��� ���&�o���i��؛��H��2���u���
��~���k}n��䘟��_x*��:��P����]�/y���or���}�!��yZ����F������A�[X�t�.����ް�'-	L�ʕ�V���eW�S}� ��nrY�\�FriL�[PDd3��?i�v@�ԁ�i�d��㫨5"��Z��~\��O|k"�1ҭ�� �7O�F�b��%5d�߹�j�B�'=&�gG��/6�q��SG8�줝�O��sH����W^��U����
3�1R_��%��i�j�&z[O�0���wt�����DT�}wf��ع�,��GjV��O('�O�-���"��#M��Y��9�VĊ�mhA�!'����3@���g��O���a�����D w�JpܕEt1)q�I�I�D��Ϭ)�:�\=���*�{d���j,�#��y�tm(�-�H<��t��~��?�:ׂ%��(���{�1F��@�@)�"p���%]
�/���O`�D��\V�h�x�xq�1�EZ+C~#�!7&g�/���qhܯ�l�G�-ĚC���r�o�.wu�rOq��>$��ڪ|2ѧr;?�u����Ee~8S[�#�n6�n�rB��17�Q��Fk))�(�,i��[0����;�-W��^��9ʲ �I��T�e�4=�`���q�P����.�m\���l�ai7���0r2�\y���j�E��X�-o��	�{�X}��b�qq�������_��t�k�~�x��4!����]P�G3�y%�Q4�	_y�,��!rn�����H!TJ��Aq喑��DϹ����N����Į��C�q��WC!M׉��"���ȷ��l1�|�}S�4��?Ҫ	�B���ݙ�J#�L�#�C0���4hu-k�M}B��ʎ]S�d����s��?��>XA��b���
3�`�t�H"�����D���/�O���A���~�Y�"r���� 6�栬)Cp-��p��� ����J��=ꬳs��d�^t��f�����H�bT�2�g���g���K�u��	�@ƍQD��BO�F�n����_hk�3�7��Յ#];��ȏ��#�<6E��K�J	g��3R��j�SJ����[�2���K>�J�?X�?�^�y�_��.��4t��h{��{G�����j: ���yRS5ݳ�	K+D̜o����))�2Hw�)`~�9��`ã�!0�����	�������@+(i��0Y@�7��1��;����"���>�D<�X�y�~�8��*��>�\��?G떭����Ԏ"(���(�*?�����|��ÎXfK^ �;�&�s�Jș��o9C�a�՛)�xh/��Yp�@�M�u�k���J\VD/�!��b,��b�W�9��@џo��+�$�/����y|����$��g	F���ڴ ����u=L�g)��I��sB�>:�1S�{�9Tr_d�`"�)�6�,���n�׌R�Z�>H�,~4���6S�S���*�)c,��딜"]���
�R�e�7 b�g��.��)��E��C#6
�����p��e )���f�ia�4�D���'L�@��)���bX�����e$�d�4B��r��.��i�����
��axB
�y�3��ʒx�}�/D��t��3�:��)��pך���A}_��5X��D��Ķ�	!�Y܍�i쌍G��½a���)��V�XD(���R�ŵ�*�q��)7�-�>e�&R�����O-�F��{KctL���Q�#�~���5
�Mf l_۠"�vw �HGpO��An��]�ۗS�j�(H���o|���!�T�B�G��}Ǖ��~��[q�D�����g�dy(��N����|�����	�o�Wq��N�A2oG�8AkK�r�LT���}�N�0�efT��^!��\��Q]=�I�GR#f��n�vs�[6ҵ>ˣ7�0zC^
,�]�y�Ŝ��V�������� �s/���K�Meش��[�cH�dì���ql͐ƭ���ӟ��u��4��D�Dj&��
�ɿAVb+�N�t�;�R���b�H��T���t��i��츨.0�f0�n��{��[�+D�i��8Ț��2`E��[����zh��~���-�KǺ����wg����{��?<��XK�h����U��V�=������Q�'�"�#��d�t�Е9I7铞���f��:����?'���O����s�eQzr�`SQ}L��-0+��4�=i�ǋ��g�=� J�R`U���pg��12$��� C=o��փ��|t�R�����	�T��U� -
nnK̯����𳪄��g��#u��[=���	@+ǌ��ڿ�������/������+m3��O/�}�������~�'cw���RI-t���>���'����.1XyY�QC�w@��QY�54���Ux��3�^���愳��������K~r;�ߤ�����0/�(~t8�y(����P�*�_J���g�^ICo�|o�lF�As�dɺ>�NW�A����� ���;�t�_�炵2 �.e�� �U^6@�ˤc?�Q+��w��~l?�Q����Ix9��.��B�;STCe��R��;V�V�|	�ف�o��:w�����y0�
XD]�V �z�,�����'�!-�J9p:l�y��1WZ��<Z�C/��q�	���'.d�`�1�!�k������[VJ~"�"=����~>�%/7�Q?�5+�4�g_��~u	W
H�Ѻ/r�#�O�	j!�e)b��uZD��d�UY��t~P&�g�8j���J���qs�H�]��0��ų?�-V�V�;�qsَ�,¿V���!C��cLR�6�j*s��P�� '�����i\�S���2�5����Gvʓ��	y���'��W$
<���i�� FXu���})V9_�����G��ᚢ<?���q���QG����^���$P��b�}�g�CfqJ)�|@�����j���}�5���!LǛ5��<�F�H){��
E�)��!�Ը�Ϳ��jq,tqiQ<'f�K6������~!5K���۠)eo�DJ?>�����v�K��V+���كFY���'O�-�
�̓f����M��&���k,�㹴~�)��X�	Am�k;�7�x�q��߹O�����Z��D�RT�q����Ԩko�V�p2v�uFxzC�c=sg�����0:�th/@��?�P���~H&�b��'�
L��+�bn20"m�(��vm�YGc�s{Xիi	:��3EJ#3�Ô�q�?��+���
�)u{{���d�f޽������v���<����(k�
�	R�9������d(��>�	u�pC��֟}zc�S+7AG�sh��SF���hi[��N9Ҥ�C~�|9Gq�8��t5)�_97{�^5���?��PD(��-Q����P䣻O�� �*]Q!*�_����2ا[��&��	���y
���+c�����#ˮB5w��?7�g�Q;�6��/L�W�?Jڌ+�6�����;���1-�}܇A���<Fc�.Έ;B+C�[X��G�Iƒ����߱�W�}�ꭱ�֡o�Ngt`4'?U݂Z�%�h`6P��;�y�����j�%C�%|v�ӷ�KD�'-c	�H�����r�uT3I��l��\˿��˕/�:w9���D�j���w�DV�$(R��Qv�ݦDwS��@TZ���6A3Ο��%�_�U�Mmt�Y:�pxކ����e�.A��z�8d��X6��?�τ�$��*?Pl�A���Do�:��v5��k��AXD�H9QIMj��V	�@`M�&�y�\n����Ǩ��4J�q +�v[�� >�*�ĺ})��W��g0{"~ӓ�I�'�D���M�̌s�Q3��禽�#�8���X�����o�֖��ۆ���ޑ�P_���B����Q@�8�����w�X�i<$Fi���i
��O<^�^��|~o�br�M����� :��7$um��vw���=�o�%���A<�f[g�%3�5�X^ް��^�	A%W�/�F WB��� ��1���D���l�K:�m���	:��I�D��(�
 *���KsH;���+�ܜ��j��!����Ȗ��"�Fp��x���*+���j(	f�9��{i!�4)�}x�2�9|,�o�$(�xӥy��Y �Z�I���Qg�b�� �ö���Eb����_��jI$HQ��Y2>�
Nf���-4��!���<��ei����1Ѣ#�������P	��0�S��S:�*H|]���1����%���'���V^��1ѣ���@Ϟ�`k8qlz�2lu7��g��F�i� mU�tS�K�oQ7���7����8kɊʾ�d��;�lp �rOh��5��<
����$MA)��bUYD�4�f譹��󂲛���y�d�F3��yװk��2����e�&���{���<(+�0r��h�R��(3H +�L��ڜ�щcG���h'�5�X��+��J�G�N�+D ���|�P@�h���w&��	K���w��NDr�N�CR9?{�	$�M�wV�E2%�l;��D����h����(J'ǻ ��]_�v5Bzw�>a&ND��"$}y��w��S����˲[��LzeO� 6�v���X�S��6�͘�T�y�����ɧ�%lU�rtj�����7���z]d8\�ğ6��%W���>.� L�À��N�Ԏ�m�$�K�-��������Z���Y�1 ^��2����}�NU� �����
#|6��MH2�6���c�!��@ں���5��	M�דV��UU�n�уX$(ա�� �"Un;����@�D0�=E ��x���u��h"����9e��Ao[FDɭ� ��ԃ3-�i�����?3]�'`�?W7�EGh��5d�g@{b)G&���=ld�&H��\�$?l,Ѝ��g*��~�d��Ͱ��n���D�d�j�C�����Y<�ي�R�ǊK�,��<?���6X�&���p>*�F�zP ���F��l��ӂ ���s��I�����:�f	7��_z��։��B��]� ��%��Ȁ�ɤ��#�?U�z��T���"���}�}�dڛ���&���\T���V��]�=�[qynIr̬k�v�W��{A��ڥRvʌ���QE����:�#ʛeWf�=x(l�G>P�0C�S�sT~z�h��L��>�4��Ō��a i�\6ܔ���R�8�Zp���D�R{�]HUز�[
v5�UN{��↖��|����o����Y�
X�{����4�v��34G�Œ:�c����ECSO��5�D�ky�!9z��g��#l�m�8�<!�J����%�� ���]UcBz|f���R�r��Eځ,v])�wq)r�n���7� DI��^	OI^Q�����̩\�$�?��Іr�����Ajb@:�q�
����D�o�y��k����]M�hs�u:��Ѩ-����84EG�:�(� ۟M O7�.Ķ|�AV����dN0����(H��AM�_�T�p���,��ʚ�F�g�.s,I�+[�$z���$՝B�6 ���e{kYl��m)Ā����`lW~V<C�ft����rK}ʚe�w�/�䔨�:�Oe*v�tB���J�'��D�N W>y��/�v-[=Kˌ��1��h�,�H8�5a�{�㉃��ui;z��]g�JV���,�ؙ�)���t��O���VT2s�e�/�d�Y�+��_D��ՠ�ۄ!�x�O����5�P���Ð�lU��:f
��FzjL�vθ?�nQ��y���й����d��>I�%�a~'�D����[��hX�JL�<� �k=��5$���,AQ���=w-=B��H��Vn �9w�{�ߚ3oo�����(7�s���*p��|��pF�X�~�;�^M�x���a�9������#��ܦ@Ղ1
��j��:���#�8��9�)z�M��)b��.�.�\��׺#8�Dd�ӟn)��!���\�-���dzh�j�Kc�e�2c�P�D��� �&�2!�BͮC��!�x�wd_
sx?�����c8�_D!	�r7�s�螀"M���3�/�7���U��3t�JO��x���N��J���ڭ�6,M���c�'�������Q��.O�G�a�Qu�zC8��{���6I��X͇�!�d�Qnu��� ���F��R!K�y����x�ch�:��%����"�ͧ��]�5�����l �iAgNGC��P��Xo�-,�%��H:��H�����s��~$a�,�H($��h�����	=��ËY�����uJc�4��`���dS3N0�׿q�\+��)t|]�`�����+�SN�qy��OP�j%��
�m�"'�e��á�`8�?�O��jy��9F�>��(Tҧ�! $�ܭ ��d���)I��fI$���^�B�� 9}c�mXb�/Ғ!��"'���*zSEUɄ� ��qƃ�4���i�]#�@\�=�g�G��˫b�� t2�/+K���P�3t���-�g�d��U)��tQ��[���q�ϱ����pT8���G=G�h���4�A�l�/�foc�J�L�`#pQ���̆/�+�(d^Sf�>�yY�R��A���G��'�Vw(�-&�j<Sұ���*˟�DO��V�g��'�bb��gj���r���vW

*���/<qf�y�E��3s��{: %�[yMj�V-�q7"������g��#�^_G\�����(K��(<�l���=�Qԋ���k��� (���W���J����d��p����rk~�'�ZLq�"F>;Q��oip��^�B�ke](ɥ��m���q�?���4�E�
N�d�4xO����U/'����>� �	}�Y�\�;"���k���?F�kw�K�1O�5�~LxK�D��f�C�&V�[ \�0�\���9'3�� �~kT���6��@�Pɤ}�8:�	�jB����4d�4i_�ՍGR���I�����޺A�}� ��&���+��`�m��-�>������h���8�b4t1Ǻ�1����i��l������4z��vf���d*�J�Ò�e;��vV%�U4��M06ԡ���hUϤ��K|��V6���{;o��EQ��g�a��d�Z��Q��Շ�z��XW�-XN?8}ϻ���7~S� 捯:;
ڰ���e83��Ϋ�ټ	�X����Ø������E�*̚��wl��_���Dg�iy� ��t����{@�����/��!bu��9���yeG,ך��B����Ǜ��na�1�X'�o����b	���}�~�B��1{��R���D�=�i|8�x(��˹�D�H��%�A.n�x䦨k���3����o���8�t�Xg��u��=4K��j3N��M� Ȓ�L��v��O� 
�A���`P���>[� �DSk�#d�I�F*~2lVd��,rn�R"b�"}]����/n�[�2O����.Iy=2y��Z�@u���SG]4�m�D��Z!�xġ ڥ��
�:&]�]�<4O��i����!$au�|��A���ݘz�0�uz�@�4��1�1/2~Z�*�U��ؒ��a��w���AS��N���]I�EY��6�fz��%����^�%�ؾ��_�+K�A��vV=u��Y8I�[�$���F�	L�,P�Q��������i��)�r�4"#���	���$t�+�\��
̍���P�b	J'����G��p���Qk("�fzB��?C��Ol��`н��Tz���ip�9�A�\&�=:���Zړ8B�Ω���R��@�H۞�=��N���8k�R���S��a���3���F)��+n�um��@W���ɒ.;2�L2��qi3M����b��b1��E:���a{x�X�+�"Ș���\_R��(��^���B4��1������CU�*� �^0x����޷o�X{�Y�!��]�'�W��Ϳ�:������[]�S�y6e:�Ĕ=I�}JBc3���s�d��\S��O�䥗�bT�G:78*�sC����c��̞�A^�/f��V( ��w@ޣ���0�f��F�$�@ s���ї���bx�ܜ7�m8�^��Bw�q�1�4dc�%	�������3Q�9]���{�[��p	S�2��$�}������r`�i�,�|"� ��]6Z��:M�k�Z�񯿐#�@̌b��9�j���0�w@��J(=����dV,{h�e�橎^(\��>�k���B���.�[D�:�*9(�|�T����9�7���\�L_��;����蝸z$m��s��U���W&�#�Ab*����iv,!���.���:^8ojV]�޶���1��l��qpH�����J��_~�6�R�Z��b6�9���jF����M|R�JKG����I8(n�Q�^��5;/�!��b���Lz��1<| ���:h�K�ĔG¾)��3w3�ż����58|I=�'���y�C\�Ձ$/a��֭p^���܃�E��L�C$/��ؠ�_Q����93�S�#e8$��H�E�a����z5y���&aj������_�XƆ��Gr3&�F�3�nkL�![7<����%j�s�C:)�l�r��h\V�IB�(1VbiP�eF��?�&�B�����:�]7���j�(i�4|�x�N$����W�B*���2���o+���6�_0�v�0XxH�2>�(] �Zlp9�aN�2���:rP�p���m�F�}x�<#�}�q�X�l���zBr`v��PS�N�E8<�cm?�ظ�{|x~�9X�D�k�B������&�I�[@c���#+�z��j�ވ�9N_��b|����Г(ů�DK��n5�swVfKM}T��dM��1�Ɓ4t���S_�@�AODia�٣�b?�W�\k��v�F�uQ{��#��{�ɹ�j��T,���R�ղMB�%�%�)�s�������P�ʿ;��ă�?S�Rz~������> T��UFn�Z�-���}E�s�rk�|Y�����f���MN��jSH�Nb̰�O�,����8 ��%�*�`�v�ޱ�3���$oR���1��p��!Yr�k�]"��UN˥�#B)rۏ/�%�
8����nE݋�=FD��R7aS7qy_��p����'��7N�ۻ/uP�����S������8�-
�1�i�ijP��kYK�97��ɴ�Ev?K�H�,ZZ��Yc��ԼQ� �����a��1" ҚD,�<��� ���^��
2���RX:G��֮�y��s�#�'>=r����*?��tb�o<�!G|V�yS����W��s��W �(I:{��Pb>����n�6�Z�q5���#%ɫ���r�=��~��'V�
l=�H�0�K'��StT*�y�
�
�ɞ�4��{�	���<۝;� ��Vp�h0���ua�э�.��)m	A��q�޺�4��U�����yGQ��{;����~Vt��W��7�yvy�X��OG��ܟp���Z�,Y������D��CH��FR��%,oY	��\�������1�t���h�P�Wh�U�?��7�)o�'���5aG�9U F{?��:n�o�%�ÜV�ta�IF�Mi@�_�nǍj5��?�3��S���|�zh�!�[�Չ��Cgu��P���յ�)���Eɰ<�M����;[���賄�b��Ƿ�P���P��b��iSU@V�R�B�`�fu[�w�s�
J�;�-�\�%�����B��K7y���y�B��e�|�/0߭����=`��o
+� I��RU2�Zv��fcR�@ۡ'ܮ��J�1��Y�np��4M��H�y�@�w���P���9.�s����&{�op k5L7k�!S�r�����G�����L�+�L7���p�~D��_�LF̏�w����p���X�.}nJ>�juH@�,�j�"��x���l���X=��JXܮy�+���g?��9}v�l{�@�n�
�a����!����
[�P��f;#s���D��L�R���&�b��B�QJ��ۑ9D�A��,y�睜��]s�	�'��SQ�qlE^m��ַ��F��i�4ȅ �V���NJ�����
Mu�{?�n��e�?�`���?�]��q_�E�`޺&��]D�³����MN�+��������=��\f^��p(���DV{�)�K܃���x�y��x�?�vE�5k��p��
�����:�Z.���,�`2�����꽏3�}��.�r��P{O��X�~ҧ�\R(��'���N�s{�U�i���q)���8�p,�� �2ŉO�6q�FH�wll����џk\?5�П�(�T0�[����qI�#3S<*�Jǿ�zm�1$�>���ǲ�h*/��_��]7�wj�L����Ηw�B���łI����`���eY��S~�3 x���c�0�:��z�ZZ��2�F�}�^p�h8���H��ҏ.�!������zת�1��W�5:�@��*���#=._�^	t������J�{�Fu���E���Gm�N�oI���J�8�1���e~�omk[������v��6�%}�k|��\*���*��?ơ�~�������6�Tᆪo7���sH�bZ>۽���k�j>i��ֻD����m�C����j������}����`�V!��Ƹ�U��B�i�������x�:����2�Y}�K]��j?Ċ�8ٌ�<>�4O����C� H�L�#��z�Z�4��&�ֿ�u]�/��c�L�?̢7�8x`�:�HV-jn*��\��Sj��dn�ȃ�ߛYWe#�'X�F����Nc �O���-"	�k���-��ی�=kִ<Gʷ�*׬FN�P7H9���<�Ul�$hii<��QBm����B$J���vC.4��r	�ٺ���h�"~'5�k����W�E��k
�c�a�aKێ�!!��tsg������WM��9JIOiϩ�/��[��u��+P?ީ�G��>g�r�Aw�(C:�����_����h�J,&�NAa=D��������>$��'+,���4[a	?0���q�/�SQ�D����$C�&	9R9E#*zg�='��U}Ğ�C]���3?�@�UN1�,�n.(㣸�'��Wks kB&]��л�쿢>�[� mnx�.܊�q��sS_�V9g��_�:�H�ʹ��$����%���Td��u7��b�@C���-D��D�!Y�ԥfv�KkV�7��k����TL����T(�H�{�uq��n�K�K�5V.��[�1I��~�`Y5�Dn�'|�8���5�7��~���O�Sm(�)�Q�W�g9��V�]�����%��+�32ѴK�_lat���p�Nv�{?Ӳ>$�B�/�����
�A+�H9$�M7��L-V�K�f���~�gۜ�� Mw֎
3'��^���"^E_��7�U������
�����y:��(�^S��|6%LJu��F�0��Y�XR�r�����s
��%�K�����)�ͫ���U&F�a.f�WP���?j�nZ�n�7J�����ƋO���+��"����{t0CF����܆8�X�?�R����R�n�9�/��U9�Ei�Mɱ�͖�B��\�(�z�>�Y5�ڭ��?i^����o1�P��迋bb2

����Ov窝6Sv؟�}��Z����e�_#p(��{��T'����xs-��}�q���ցm�{��j���r#�1~�<�ҵyPi��`��;Q}P�aا��ߚg�䡌b�w�&��2��c]F�p��D�!0'jR+$�O\�-B�?��;�oAP�%6��f�.^/G��ׁ���"q?��+|���ѱ��⁥����o|y0_������cϻ�dI��?w�K����������d��o�M�7|�8��}���"ɻ��գ{��$�C�j@+~Yl�N��ԫ��^VZ�܆Q���a�~�%��b�ꂩv\~[4J�����ce~U2Qw��dA�����\Y��,��-NN^������>�<� �5�+��"{�2�,}tN���FW�ѭT�Ɔt0QU���]/ЗbQ�UG,8��.��[�݅P�q��2���1�}�n�*٘_5s{���d�%��S����}���4��h�/��n\��(�
A�~��k�{5%��Y
�(4E���
]�Ӫj3����sń�s��v��6�9F-�"�3
8���48���B��T%�P�6a�Mk-�^�;���<sM��Ҧ��\�٩&">�5��3����9�@��r��eM���T_?2�+%��\�^s�o�E��RX���*[2%s��Ɖ�YKPuw�q���q���	�9R�N�.���x�-E�o��H�f��XM�����6��p��9�;���
?�T:�)w���t�D�_����n$��ǷU�f�ݧ�M��^K��Ya�S��������0��<�0�9��4�F�=7��v���3̝�kj��f�;�\���Z~4��5țRkqT�ֈ���I����ސ`m�gr'�5h6����)Z���(����IM�^�I��t ��dy^.��uq�+7B��k�m�iv��P�ˎ��דCл`����z0gLo<u�r\�rM�b�D������+X@�$�c�I��(5#/�!�˱�I��P)��
R��{GBw �ﾽ���&L�����`���P�:�M)��&0O�O�L���xc�,D�=�5����5��̷��|yaS1��M}M�fE܄�q���-)�LN'���d��8~j�Zd�%E��g�0D�A��I1�OӮ���l����%�)Z�MغE�#_=���h�X&פ�H��#s�Gy�DI�侤9'��-�-۸�:Pu*B ���&^�i����sx�n�x�a����=N_�n�o�5X�cdg�g\���R�!��st�H��b��l��Ҷ�eȹ�C�[���)l%�;��2Fd^�t{Xd����M�X���
������\n��i&�<,�VC�m�X��3>��#�TR���?���B[���*�$n�R��?���<P��H�����m�5�KV�Q$x�u��i�D��p�7I��W��.vX��#�������E����<���Z��a>)�\��w�_k�1��pޓ@��A�h�"�w�725ڍc�YM.wqo9��m��.��&^� n�
	�XS��[rT�Ѓ��ƀPi-��,h;�6��2�2���*ϰ=��v+�-ۭ@Q�Y�:��U�r� UC��ans��4
ϼQ!��#�V�a�0�֘���RX���hy�ğ���B�C;����Km���Zl�ذ=b��q(mA����Ʈ��u����4hˇ�+����D�5ŧ� l� ���h��!-҄�|*��f�9�����e�_��Y��\R�?h`gܦ���Z���{�6�p��p��:��T�HR�_s1>��_�Wh�z�������,�I��S�IFK\���)�B��;Uw ͔��h�3�7!Q��(�wuL=�D�3=���.ޔ9U�ce�����T{b��P�zn�D��dh��GF?X�ϱ�:�,O¾ ����7<��Ր��s��GY>v�;p�6�sH�FQ=��\�]y�9�aa���M����b�=z�<�@�Ē3��؋J��Q���в����?�]Tj�s��K����Y����'��w�x���~�ZtX�^��(�9�
;%�/WT�Ĳll���V��a�N$_�%�ZWkfn�#���m���7��OҲ�iO����XKY��[�7�oX"|�h�ё^珛y�N�c' �=���ls��E�"я�P��-i�^�.�#�V�W�V�-����N��?�.�y��@]�ӒZ�-�}�@'CRܼi�!s7�X�)�2	&�ۜ�T	%��6��I���ֺ�s(2tDZ�_�q�Ʌ$d��UwIn�hx���������Ȋ|R;�.[`w����Ybj��P��� ��z�~`ؼ�i�F�b炭(V���]o�;�ۄ�>���%��<tk���~�]�!1rSv��l�UN���9����խ���S�y������	���1�;����:tլ���ZJ�����v�@`��=fA�>}tLq�,�D��[�U�IK1�L�������d'�3e��E�T�2P2z�������?���/�}2�y�UU4�T��Q�T-R�ނ?G������i��#GB���=�AR,��<is^��j���p��`��nS;)�4���``]�OQ�R5�Gʮ�P�>a�\���uO{���ΎO2@�᎓4��@�!�l��p}<�zV4o޺�~�GN���U�Q� ������Uu�=�w�P
�{8ш�J�J��I���ـ&`��i�˪&��s�%�� ��\3��K�_,L��7���iG�E*�%3gѰ�Ҍ�wr�͊��Ӹ��������*$8b'�a[�mvS�[R/b�6�%�(#eٔ<�A��L��4�?!���<��I���.��>��ob�[|��f��j�G���$�O���ɚr�zd)斪�,<ݬzP���{&� ^�28騬�7V�\��bW��2y3VW�����~w�+r*�:��c�7iZ��S6������*&.'��[�>0�=�T0L����i�	����"�����(�ty] S	��aC��yxH2�K�Ҟ�M6�:Ԣ1bt��w���!�P�h��t%�Sm�c1��L���y�+��j��ۗ<b�,n�}}I�S�d���|��d�ھu��	g���
��SN�3N�U;��e�On��O^���c8��"xj5@�
gb����Up�=�o�bk��@����"c�B�#��w7aV1��m�C������Um|e;��K�^�B��Ԙ���'� ���m��lUc�dӸ�~��}���-����f�4\��5�DoUW�	����)�'/�_��Y���1\�Qr�v�[ݬ�]���}��~�]��GM��|vW@zr�� a��/���=�B_}\�����QJ}��L�5��B��
�U)$V'&�m�I����r8�|�CNv/Y..[�Г����^*���'oV����%{rJ��xH#��Q8��{�uk����sR�2r�ýr��6����^���m�e������ h/, ���� ���$�}���R
�h������/�����k��ƛ<Q���N�>��~y�6[=˶�K<5)0�ƌ "��	<:f�h����u'�F�֎�r=nm��w�|3C��.u�k���;z+�lʏz�#u�r5���&���D	�6�<\��!�ˎ.��ѐ��%�n�na�MB%���k����QVN,[�F�Vi�u>8X�m�z(·gj$lWdyj����R!^�`��a)hĦ��+����`_��E�
A^,�����`C�������w��~��J�gD�'J�ࢃ��<�l�L&���ٜ���b��^�4�m��*�T8W�����*����4ja^O	4���=B>�[�͜6����XѡK#$X�yI%��ۂ��+��
T�ړ�zU9[LY}L�Dd�c�׳3B���fNWh�Ur���du-P�x��;���9&|�fp$�3)�OW�	��*���Z��!�S%!,&�^�MW����.��!1���@��n�$�߬��� ��F���|�ߜ���QU�C${>����9K��l��tq@Z��x��q}�z��o���?R�;o����P%/�4xm�6֌�S�̗ �'V��M($��Ƨ*hx�_~��=�Y�Lﬔ�#kZ�-8ca|��[���af\�'��~q�̐�߫�{5ӷ3�K	B���H���	m�â;�6|(/�h�1�~�*��`�'�={q�y�|7��O �����Ж�Imv�D���{��B`yHZ�m�ݭ569���A��s���E�*e�A�[ՏA��F�=�a���h+e��`"&��,���]�`��u��:��%�og �$�)�$�����w���(�jwJ+�~�&���J�-��B�	i���_9��!)ѵ�~s��`m�}f���T�pڎB��7��^��Y�,��� ��@>�Rr�1\���R_&���$k�VO� �E�Pa��R����@�C�5�#�%�n�.B�un��s�����#�L���!�ܖ}���y�c�� X�T�Y~��W��kqIv���4)�Q���H0fe�5+�*�(s��K��f�,?���[�����Fɺw�?U�ǧ��塲���R3]'d�C�u�Y �����_��Ӎ};H�����	_�����ڮ	A�E��U���|仮�����rbf1=O�g.>
E�\J����P�๓�a"#�`�2Q��a��,��;ҾO��(�s�u�;���M�FA?�TjR��h�R+���Q�35]ԟR�e�k9�풠SY�DF����Ճ�l�IA�>�?�1��׀�J}J 2��w�Q̷��F_'��e��{��g5�bf6[.�D�]�/Z��n�5p��6^vz��I�F/=To=,uڄ=K�����g+�0r�1֜�;�/v�O֜kN@F�������4�Ը���\�m����JJ�c��]�d$X3N�ެ^$`���hD���w���b���z�u�ԅ?3?@ [;ȥ�vj[�o^���k�e������Z�ȲP��Y�^9)�O0)�l����A�r֕a�#�x`�i4&�-*���T��������k,1ز$��ǄW|+7ha�!��KH�H$E��}8�w��3�@��y�Lڲ}���K��L�'�S����-�$�AF_.[	��*n#
3�unW�M�UÈ��#m�x��P�R9^�fyh�0!�ݢ<������Q�bՋ�r 5�EGy��Ϗ�;�i���H���a��9�Y�y�U�Oï�q�Φ��k;'n�:�!0�_|~>���cNd�f�j�k�d �}��j͗�~�9���(	����&�]�j�E���LD3	�x�E�F���m�����0���mڂT��7��7��,ZUޠ���[_�릅�R�@XW?o��-LV�#���C�H�ˈh�(h���𛻝����}�и�<9
�
��cÁL|����&��MT0��������jMv�Y~�g�^��RS|�����)a}��h��sJ���f����r65F݀�L=��WX����PUK�����l<�9�Ǒ4ٞ5d�̯	�"!:2K�Ce��~���H��G�*-�Ne:��Uv��+b���t0PM!�L��+�'���+��X�E{ݹ�ۈ�Jc� ����ԄqP�C��;δJ�X.\��tZ�F�1��:L�+S�Ujk�~%��G���L��,��Ɯƫ]��Y��>\W �6Ԗ��.�X.W풛��K�d0B�A��gZ��T�������ٟ{��jR���3J�!�]��ףZ������C_kt�Z���+�z�`|����#��4��ܐ��:u�?����Y��{�|t��r�+��S���_�YV��q�i8�����O�#'q#�>�y�������mj�i����U�s@?.M���{��(�2�W�%.`�lK��~��Qߏ�-�W��;ʲ1b���F?^���])B
}k�l~�{�)C�6��M`>��XY��e3�4z��_�,ș7ge|��\����u��Zߪu����9�|����3c}Rж�h�S�S�t��u�.(���إ�O7<fQ��2D~�h�[w��]�ê�8����h�W�5�ET�n�$)�t�J��<��ꚼj��nS!o�N��
�YX�z���G<�9��pjlv�E����{�#���B������u�#�ղ��/���&Fp )���k���k���`��d6�!�9�O�>�2 d
�#����T�����o�u���%l���*w9�����6\����O~=�9(R%��HjP�n�uƟ�째��P�X�?F��T�IF�\BmP'1mWY4�@��N�N�!ʋ��>�k�/��I�h�;f�0�	�G���8\%�F�� ��G���u���n��Z~�)���_��'�����AzV��x�;6��jm�	ݚIQ���@P&��kw���=���-��X���1�v��䭿�y�P�Knqc��V� �� \��XX5q �-��3��(S���4=}Z?���f��r(~��]SR� �����
��]
���1R�R	�[^�D����X���u��F��2���T�$+%�C��mﰀE��+��<�"W�w�_%.e���&-vf�0���>���Pѐò4�ֲ6����^?�
���|��,�,O�}�u���0j����`�$���m����G]Ih1��]�yN]ɋ��'8��xբ���;��*��r������3��z�s$j(��`a5�%� ��5Bo��	Y7W�s�k�E�lA�p�N7���a�>hzY@e˲�Fر�&#U1�-NM	L��Q � 2)Q���p~�L4H\�+q�[n��G�Ȣ��s/�T���U�c��{�S�����7�P<PT�5G����/Ti0��X��q�ݤ>R�ZjQ��P���Q���Jm��Z)}�U>c�b��fW��G0����/��Dp��k�U���̈́ű����z��=a|�Pj��$���,kƵX"eB��H�_�� i����ǲ�eR�-����^u�����l�R�OM�e�o�0�	���/|e�0C~�D�DJ�
�L�+�}C`�CNkb�������W���nS���|�'i�6T�f�. �gU�eV�J���E��i0$�D)����K���XX\���P���!�eg^�V"`���|A�� �u�l��R�_�=�sklYdqS'���E����^v��a��\�W��ټk����>VwF�g�00�IxŤU󳗅�v�x�ʹȐ�#�<��q�!��Y+��lgbg~뚴
��KKq�zv��1�=��1���õ�3km��y짃�F�m���r"���W�������G��Қ�xx��U}yg��YA�C��g��B<
�ſ �ΆwO��2hӝ�i����L�5��hy�F,���L��'h<�Ƶ�"���_D�6<۰\#�P�%{<��<x�nW��o�M��f�ޅ}��_�_W�hLʶM7D�
���x�m��,�ռ����X��$W�`nC鸇�I�b���.5���`�][��w�|}�?M��v.����G}r�B/=�7���q�*뽪N��2�؊KV9\ci�/��a�h��+)�ˇ=�S=+���Fw��W��Ҟ�I���[����f ��'dDO`�̞Z�Ȋ��by�ƐZC�:RCC �v�@`88#��`P��ydr��C�#���ɛԘ���}�֬�PkLҺ�X��pb����hߧ�[�R�W������/*�l��cd�I���"����0N��}�ɩ�XO�,�C�C�S0˰�м(��Uɂ{qD�_P���8}(��K�Ku�'��'�>��&iu���7�i;`Os��s���W�5�}�D�+x��O_�����)�:9�B���0�O���-L�s�.� ��@���:2�B��`��=Z+���
c��˸���.��چ%h4�Hv,躨M=G.�HβZ��'v����q��B��\���G�i����"\�Y\/	��h�k��-�R=`^Z�k���Bx�)�cޏ���T�6��M7�M��)���>R>�D=��7>_ZБ[���(f�<��k"gp^�Q0wQV�~����y��p6���V-+�k�з\�^�u.�����yE7?�?�e����Q����2���#��ҫ��*�½��vT�{U��bN)����zb��Q�q�5�p���̪����Bc8��"��h��ͱ��,1F��o
�b����%3X��-Ŷ8
;�TXUU�x��)7p�G�a�pf	8S�(;07Э�5�JQK1�����3�Sp<*��V2I�Pl�d���u<Gz�pm7�꜀��E���rM5���N�bmog�C`
�lb��}v}� �"�����A�O7���:�H ��>��g�ɏNW�p��2�ɢ����^%X��G��}:^b�ލ)��I+���G�KMG ғ-vEt����k-�Vֵc��ݻHqfN�D������f~���U���:���5��+_�g]Z~�9w�,�/��_�ג�˩�魙5j�Hpq��ϋbq�c:A��	(��yl4�`�}�\0��}i�g@>xo�\P-����ŏ�������3�q��Rޏ��(dlCqn�0+Z���
\�2��񤋗_�P�m
�GD=%�d�,����NƂ�E�
?&�mFa�I�&��1Bd�@�	1+��og���= �{�i?����
0���~��E��
v�:"N�,�x�@�6���Q엒�˂7�$�u�l@yIL���E�y��,}�j��x��������12������V$p�b�n;cT,`(�>�T�R�3�s�zo-۾�9�ш�<�D:h�Zj��F
�n�ڔ�؀�)���Η�F&��`\X*t�J��I4�q�!B����h��^�V��G#�7��)L�,��F�(q��w��~nX*�o����kcA�o����	LG+FMؘ�]l�`ѷ�P4�X˙�k��_�8���MA̰Tk}z���P���c�����g��& s���^O,/�\̗�!Vx��X�D�{q13�ʆo���L�����-��`bp��R��U=f�&�y�q�r�/� t\������oq�O7�k���r�vV�A^ ��Ҝ���-�8��g#����8��i�3��#{�L�(`A� ��ze_r6L#�X�*�Z)`���fg4?���,�6f�P�^%�`k�I��Mx�a�@76`��6硆��4W%,�v"�h��S�u�q3|���C� ]B�&b�Fl���<�~`�aĤ�c�B���}�(�}<=�x���¦�T��Soh#�%{θe��	`�xy�Ir,<q�)�z�e��'CD���߿K>�'�1U�t�0W��㞛
�C(��Μ�f�Z2p��0����gpԟʦ��-/�h��P�� �0���z�$��$�����7����<�#kG�R����2�k
I��
����)�d�b秤v~��p��Ӿ��͊��k1���`�#���%mO��*���(G6���6wp��B�� ws%�$��:�8�SD�����T!OEWoI��ktH�m~�׬����5���=��!\�s�1��>Z�׏�Q�a�J/@�MYrq�$���AV"�{��T8wi`yx*�$���6<��)7KH��H��d��jHmI��.#�PA*�Y-��
�t	�S�HՈ7�!c�х����p+a��+fWttP�9` �	��C�[3�M N8�ڹ)>a֢��E��DD|�YcHF�� ��T#Z������^`�(�M�h�^#��1�VHtс�M
�?`4/�b3���w}*��o?�i��*}�^n��4.���a�%�	��a�&�Qp�2=O�h�;%��0i���	�v��y��gn�ٗ���b�[�׭U���a����41�=Z$jն��q����+�!0ԎM��|l���e�>qcկF{Ȉ<���uJ����}�n��R�VK���Z /�nv�ZĎ*}�ο���Z϶y���3i)��K�$�oi��������^;���ާ�cqc�<#�2�q?��t�K	0dÕ[9_y�;/4(#ܳ��f�JJ�gG+uҷ3�®��tZ�5:�>���q9��ͤ�!��e�,�q���$���q�nWu���q"VMZ�"��#dнJ^��4��h*�I�.�r���-s�t��Ǡr=��=�	��ڤl��U�d�D` �c6�*(P�Ȏ#6+��N���;�=ˍ!�N+/G�t�FUX�]��@#�p4{/vJC���k|Q�BI�R����ҕ��b�|�.���P���`��1o��JGyq�*Xj{�9�j�_r��o�`䷨v�trAF�A��+ʁutD�U���Eߪ:V��d7 ����LC�p��Թ�P�{�M6!M2�`W׳{{�YW��Kn��	�TUDJ.Y�,,/�8��5a�Gk����[L���r�1�����
g����e�ms��q27��O����m{͏[��ٷgC?�WHe����I�jˡ��l�ũ<5�����Ar�c�mp�En��U]��H���h��F��cz/��u�O�8O�_��e��IIG�v�q�y�����#	��=u��Z�n�����D� B,�f�zl��)���'������&.(�2k���z�.Ӓ�7x��`�+����r��c��k�j��X�S���Z�u@��%�;z#�h��P ��_����4%F����wH�e��,�N�xOV���4�OZ��Ԝ��|P��w���0�$�P`Vd�x[�Z��^G��?�@f��bv�پ1�5Е��c��Գ���G��<�j���f�ܿM�<�z�^60��[2z�=���I5���$��c��tT>4�{�$��-v������H7�B�?�=��2U�d���Z���)$lK��;�ʆ�z;5_�
\
m�ӯ޷�W0���;�c��f����I����pd[��6���Q0�]�}��)5�������{�Vږ��/���2JL��Mo� OyRk�,���g�9�'��TF�����@�d���h���D@�����!��s�++/4�[���n2���M+�M�r�3��k�Vǆ��st´8$m�ER"ɏ���S_�7��'slm���$�i�n�YrbIL4�_�|D���l� ��%D{� q���lv�Y�����Z��[։}h�#̉MH�i�*x�i>n���R��qJ���XI�#��z_�d��>�3�������^����^JSR���)!1%�c�u�nŪ9�\j��l�[������p���&v� !֯�B>�U!u�h7�bT�u�G�r9��iEq����g���x��@m���ʛcfj���,�W�	�N�a���1pS�vj��GRF������:7��59����K8e.QjO���[,l��x�����	�FR��b�O�������� �J>�!"i�)�ݎ9��� J���[+�F����]݉�8M����["����W���HK[���Q��R��G����Ƥ`ۻ�������8�~J���̷)57]�GQ����l�v5��U�C����)�Q6��S�M̔�S�I�3�gr�p�K�m���<����W�-s�m�����٬I�LB�+�'��w�K�P7چvd�.���ӑ=��3���/�c#�e:"���T�XZ}(wxa�|؜sb0+�4�v	 >��ϕFa�����,��5��a��dr�>���'��'[1vl����@g,�<��&��ӡɹ��͙�[P�8.r@�R8��%�2C�ܭ��Y��~�aZ��,9�xF9U�A=�"��b_��%⭂�M1$~���{�����w��t �R�`�\�}��L�A9��:��H�|>�+�<8�Jp{��]��H��A�P���X�������[��
!"z�{�*0����Cq�����B�fccۃ�C�U)��T,�K����"<7��Y�05=VJ)��E[_m�0�\]-��Z�����{5����J���WH�-`��2�4Mَ���<d�u��0�a���]_����a�fY�:n�$+���:`"t}�ynbޛ���9�F��'|��\�fv3��it��%a&��A��ܝ�Q�,�6:	M���Ĭy,B�� ������1�w�m{k��mWe=���L�qݾ����6`�$�d��}�����S���� �Ńex�صi��5�N������aܸ>�ЄF�t�V��YU�k"�ؙ͍C~6��bdJ&��s�Y��1w�`�w���m�)Wh�\�CT���&�B��������m�
�ml�T�ߒ=]f�;8�W���٥�Hz#�8k݈�h�w�21��Lrz�}�f���ZߒV�$؉V�h���n����6�y�a���ָqI��7cS�{��\��@��H
���lF&��?�t���Ccj�BRܺj7����G�D���>��2w���r�Զ4��2����+�h?޲Y�h��g�E��w�"�M��h<2��a��;�<P�0���UBiϬ����ug%�n���F�E7�d#=^[��ifݮ-� ����y��ڿ��>:UW��`�	�l�>�9�<�)��ip�����c=�9/��\�
��Q:@q4Z��Ȁ1�usV�k�23 7ѣ�ȝV���д�UE{��\zc��� ��b0z��@ 	M����qv^%�wm1�YL��[��wm��e��'0+̫W`�V�sj �@t�G/ۃݵ��]<��XVhF�'��7�L�p
Nzx���u�4��x���-^(���$��k������}Dr�سˀO���/�2��B����|Pm-�qo���`� �S�.;*�0���0�����o?�D@9Q���7���6�(��Q�lPpi�;ͭ���Ί�:ߧ�r��-G�d;�V���l
���~��^!]�v�a����O��{F�.徽Q��uΞ7�I7+Z�_tT�����F˭V����=hV�K�:Ҭ���:�9�Bv�ËU=+��<Y�+�uq�cڛ�b�#��@O��5 &��,��=�K�|�UFGD�q�[�q�$�_��kXu�x����T�Z3��t�L�vKw�3;K#����@N�b����!���'7^@^����8�^�j(�O�|�Cz����8�弑A�C��m��J�����!�ċ����23ʣ���z�<��t�oV�!+���6M[3�Q�J毅/aRCT�Y���
�#r]�^�]Fi^��{8�?Pla��e��R@*�ER�L@�Q�y��1U���z�_�[�v��Ⱥ�Dm3"��� �Hw_k8�g�����ꣂ(ֺxW�����Z��K���Y������V���8����|�ɉ���W@��C|8�4��C~���R"-�8��F��E��U7	�]e�.���32:�C*������9:!Z-�2+��_��\�2���g��Nr�M{�_3�ԇZqUZ
(�N `$�yJ��?��Ae�ȃm!.d�M��k�����xԣ�GC�h<��-�UL���	�qu��#���~��̀8a�w��B��S���ݨ>D�����P�ԡ
 ҄�=Uh^NP�d\��;&�����Ƶ��W=9p'O�d��E�C���y%�k���>׭���rx�H�-�ƹ� �R2���F�:�u��9���>?h~�JW풥���������<��]4ب�6��dڰ㠋2TL�=l�(��^s��y{-b��K�eJ��1ic�z8��
�L_��`����Pw��$�bi��_R�/8y?~��
�iqm���(�vf������2���Z͓#���T	���i�%c5����d�UW �b&\�;�{��6-�������/���g2��6s�N���Pb��w��R#т�� l���Q�'��&���u��`��`��կ늹hW�R-}��Q������'�aG�m�	&�Y�Z�L��A�A&��9��%��#m ��Hq������Z(9V���	J������� 3�<Q]Yt,�f��Τ����i�ev{��F�R�+�rN�;C��\���\�˿�5h��"��P��8;&�@�@�tSc\_����eb@O�o�^����c�i�q����^�7���N���N��؜���:��vb���_.�[��`�W�4r���BN�
��;++x���S7t�6�ي�
<�'6UF4�*R�QYO��`��OX7��˼/%�Q��L�M�qGk��Rv���7�G`��B��;H&>���+��"q�"�<b�� �S�D-�ˬ�`_�T�]�{��S�O0]�ob�� ����|�eP=]q��=��cD>,��ܡ`hD��Y��w��L��������7�w+�8J�c��ꋑ�����^\��g�K�M���w�@�'�{�RU��A'[����a%�s�ﺋZ��C�r,E��D���� 	o_��'��*�#�Qć-��5���>:ɠʁ44s�d�n��B��/_��������T��8�C��cb=��	�@�E&꣢�*���yFJ�7�+�I1d/�|��J��W�~u�z���&�u|ǚ9�x}��3fJ#�4�Y�t{���\az%����ى����@��ҕ��	�sZZ���g�-9��B�Z�O��"���!���&rt(���ﬄ.�U/{�{q7�*@���z���6a^2?�!�����p�~$�l"�B�����e��sK��Jf��%��x�P�_�)7�ȘgO�Y�un�����6��8L����Ǒ��?�!Z�C�R�c9�%�+�����"�a4^��b)%d��	y�4)ܨ�r"Nǳ b�����~'�w�7�x�) y��ʉ�Z+	ǝG!#����%{W*N~&�Ùg:�g�Z�(��JQ}lb�W7�?� ��ojn�
 �|ƽ�����Shצ�,�7��C�����Y݊+0�5���~�z��õ��������	+��&�6?��|�U#�X� KEoN�{@��"�|��)-�:�d=(���u_:��H����(t}=O$�J��@�$_�sz�)�h��c�*v*ʸ�R����lD�':|�ȕq�3b��܏��	��ۍ���-��U�鯹��u�Ŋ~C�_�6F���I�嬎��}Y�B�ˬL��.; �P��t9&�خ�[N��ֳs����>3P��Y�*��u�������!�F�ߔ��;�繷�~(l,������Klp�*�NI%�1������ӦF�r��$�$���EX�ng���e��է�u�{�粸Mft��C���*C�/*"$�l�g���æ�K����qdYq�5r7�.�~,�^���"%����#Ͼ��t�}[)�WY��F�R��ݪg�V�c��뉹{��w�bS$���[�����j*�sz-��.~���CI��wP�/�WN�G"Ձ*	F����fz.b��)K��w�H�O�4�TB�i'}�s�����	)��9�[��|T�=�o"�Y䊥��w�׈�]5v�N��=Y7qӠH,�UZ4��9����'!�JϠPZ���QJ8<F�K�#����I����/�ȴ5>���c���~e�!�N
�ՓT�=�ަcP������f-z���U⨒BkI��ix�	�z�^ԒF�` 5��^tou�
$ɇA���H%*�*a� @|>�=Yn��c{��<�`M�PS�:r�u��[Bߔd������%�"�|,�k��ۯq�/�<R�L/�+�3Rw�P�4~���.|%��GJ���DF��}7Vl4ӃM�1Hq)��g�\\]N��L��,/�3�B:���K
��׹^d���s�e�Ȫ�����ѝϫV���@���ݓ��E��	�<9ύ�u��IV���!%��5�JzA����6����ǐ�{N�a�gѺ:�Y�/ A(�ͿZ��;�ioŲ|���2��v��<C9�@�GVSc��X�zʳ�1�0wϓ��_Mq���{��m,�u���N]���&j}�c#�b��X>����!�!�v�(Wq#�E�eN[�C?�F ̩J^� :��9P��ơ�+5�w���[��#9 �s`ƌ>��V��f��N�ksP)�ۂ�*q	49:��G�
{RZV�D�{��d�Zv�繣�(����D?�������O�Ԃoў��]e�e�z�\�;�+���&�(B�tܖ<2	1Q�z�_�h,��-���ܢIo�`+�q|����I� ��뉐,�����zv{G��������g���H䉅8�z��3�Rz�����"�E[�W0AV�S9G��1���(�
7sj��Ǽ��6E�#��"��8��YQ�H���@�4l 	�5p<[;X�&��W(qr=>����=� �_�僭hh����k�T���y`K����p1������W�6�͖r~ ;��߰�q���� &Ӏ��J$A�gq0k���rp�� ��g)��3��zNZ�i��ּ����`ݿ��<����x������mgq<�����9�eO���g���3��N��օ�q�;�6F?U�@��w>_I�@�)�=i�庳���0��7.�j�+����͗D�.oഗ�O_/B�1QY%SM�>��1�exo�
�6��a�ˀ&�#h���d��Q�ԑ��qN��]K�ܰ�����M�_Y���>�
����ɫ��7��[��n@`�g�����1r���Py�C	���n݆�b�m;{Ɓ�I��X�F�&�l¼�(����� P��ѻA�0�?E�W��q`"_��?�j?��8	�T�,_8c��� ޗ�0lUx"��N4��Ɯ��*��W�+,Bۻ�S[�S�V�(!�%�S�v��_]��W {D�v����q]䁳3�qP��Q�~Z\�~���'j�%��/��I<ypA�⯨��:1�N�$DQ�ȜBz 'ޞ�{ 1��ؓ86a���C�PY�t�s.���t��V���c�W�[n��B�Wq�%Z�O���(17�}f�~����� }���BKvu�phҾ$�;5�&y̖��2P���Y�mst��>/�7�)��' ��*K����H{����L^��D�wCZYVa��)9�z��Ǩ��4�ӡ�H����$�����;�	*��j�1����W�v��a*��j���5�������H��*�|��Q�7֐��jf�;s�S/���巻v<�1:�q���\գQ����3�^P�&.��@M�s]���(�	���B�:l���Ω�4uS'w+��>1�\�0�7kU؊���p?[����`A��L�[5ɣ�%��ø>���3��~v}!�}���B�DN��V�J�d���k���Ά�?؏�$6C�g]�b5Rݔ��� �iN�p�]��P.��p�;�c�X��5�M>,���y.�B�EhA�b��l�����<Fv��0�쭳�}���2��NY�[3v����?�ԓãC= ��y1�E@q�PJ�i���Op.2�&S^ѿzE)���o���vޔ���v�' ��cԑp8�$}9'J���a�*'_KN�7K���K������_�Ր+`�ѷ����9�
��y��3D-�!�����9�	:RT�%�ĉ�F��*��zh�"aEݕ`P^h���S�G�$ۛ_C�"5EOC���/��{��QTWTj8���\��������3t4	Ci�����q��I���4�Ҵ������>6$kJ�j2��w,�Cx��1�����Za����2ι�&&�a7.�9yߓ�@����,G.�f���#?]�KS�)�Q�=�p۳jk��cR��,tVV2���j�笓�����U�����[��C˿�1Ȭ�zH`C�uL'��z�
��M5���m���zv]���z-�������Fم:�����*.g����孫;�� Jg�q�A����\מVV�}�~�NI�;2M��$s0Q�s;�J ��ڳ�Ӄ��"�		TZfqo`V�vHRt��I{�+|���~y��v##
�3�S�vk�2�g�@T��<E�Z���"��%�ԨE#n�E��8�#=XƐ��i^��Q����~�y��X�W�����o���	�S�E#�����m��.Z 	"���E0�ze;6�^�N��4��\ը��0�7A��v���>A�5�^�ϰ����V��Z"�l��֍��P�J��P��mU^�c##�ejc�T�FZ$�*��m>fd֯�FY�h���b)��8�|�&�@]D0�/ g?�i�S�(����1���gC��&&N�A5&SD��1J�R��H�%�,�i�u�H��4�|Y:��f娓����$	h e�h�������b�)��`�=�w���[�(Ec-xg���
XR�'jW��B|�N�z�F��$& O�'5$�}�{;�z��}�����ڠ��Ɩ��h�A�q���ةV�)31�s=di#����A.� S���Ɪ�̪M%���{��(<S����������g�����U� ��Y�6���]\!v�l��RT��c�6fʁH�wI��Ԅ���R�SEV;E6 J�uT^���C"���?H�~�Z�����(�/]~1;��O�B�����
60�^9)� �B�¸&��Q�����`j�t֑��+:6���z`�'.l ?�H2��Ln)�D
�c͗3B�nC�ϲu�E���T���3-$�Rd�<x���i��#��9t���gpx�U+v��9�rځ��}�&��@G��ml���0�䣬� ��]n8�����l<���T:�h���ܑ�����=��۬g4PQ��E�v�1��YU�3e�Am�}����y��R%8�0�Vg�Y�El)�x��x��p ۯ)h�y� B��u�$���kqX��[G묍wÊe�߻W%���8ތ~X������2-�� ^����[x�׏�=T>[W�V���&(<��empÄ�j��R�̪%�+��(�w��;h*8h��f���Y�T��z��A����g��[��3�v�R��-	��7��4�A�����u�BQD}��6-����xO�!�Et�7R�`Yb6��ch-��*{��\yȪ�ϓ�qG��a��`��◒�`c�d�\�(�[!q6��]-��7���5^yg�[;�
�UD����p"��'��Y5g��lJ�P�A���ι2([Q�Ek�u�"̽S?�k������a�C�}�su�W� z��ۿ�Kd\3�M�੣���̌/%b�m��1�����MrTMcSt4�w���O��8Kaj�V�Ug�믡���⛂�}ş%�*�&4���9�XH�#��m6C�^�bX�����ʢ���A�U�ͲA
����=�߾��|�+�W&�ݮ��iq�����_!��84q�0Aӹ��-�l׮�7S],
<��j|��1��.#uO���p�a�w^x�(�������;tP��s������沮?�U�|����	��W��F-�ַ<�l�SP^2]��f��n���yJ$�rJ�'Ia`;[UV#ۢ`uXy]�@�4z._����y1z�;���j�Ym�o��ti���eő,�D�,6Û!�ٴ���b��eD�y��4F�B�8�ߚuMXq��/�:��<l�n��`��W!Q6�O���'�B����� 3X����t.3��D*8g�')�I�/��acF���CȈ��;ұ������A�[Sv:[,3����;!�5�Bc�����'���}Vo>�R�_�_��|����A���@��Ѣ���rt��8	��I/v�
�讆o���ݺ^��&�Pe?U׷�)�D�Q��L�	����!>��k�q �p��zs�))��ng��w?rJ�s)*��������y'�G�U���G�dG��DF�5�����L�O]3�^~q��L�ǲ������3�o`���6J�
I�[|�n�8�|����[�S����o}����04��LG U��Dm@I�)R3�6���VOx�Y�*�Nf�.JI�S�(}�U�p{�o�#�͘n�2W�5�;P���'gɑ
��n�޲��̤z���W*�a���Aq ]�+��� �@�\+l����]�8�O���QMa���y���H���z�p9�L~��b��d'��Â��&���bGb�wJz��i9�q�^��jM����#"�h��c�p�&^�9���(@ ���&� ��3�{�nw�EU�Wص�byp��9���}�����o##4n}�J�_��»G857,mO��ǂ�	���/�D��)�b�1"E�@��S@r�7�J���~Nc;��\!�F>G+�g�s|���y�_K.8	������=�ǒ��Hf��K׍�O������*#�����kٟ�m ��қWp F��������V�ӯ�yD{�l=��T;�pO��E���ά.O�q�?P��G�(p7(_X�ȩ���Ҍr��t� N���i�%"oћ+��H:.ܲC�g8�~����&�~��!��l����|�.��\�NAǧ��E�衏�A�( O���>X0ug�q�lj�bn6_�'uvL�L!w�@�����[R�o���:�$܊���s�S��c�N7���qaC�	A0�)����f�H�M4�����gD%��W-so��奢�R��L�4��E��	������h��C��)���7����@W� �R�hD ��>��A�aY(A9���<*�q���X~|�b(B,ԠO��\
'\���@E�9uĊ&8|�;��od�vf][�g�(J�v|7s�ia�#w'�]%��-@��o\��Bu��Dq��F���2��{�\���3� <���E}|�|%��w��/�Q9ڣ8��,��[058u$j�ψ�U��vՋm�1���S�x���ʯ^aO�oCQ��Bw�U�R���SC�ڶ���K3���;��t����4æN/��9����w���v2JL��d�� ����j��%v�%:k��z�X��Br\/��f~@���K��+�͹��D%�@�7ȧ���-$3Ҿ���Un�9M\S�ل�9 Û�(��2��H�z�E6�"̦{�5�=�6q	����H=
"���}3����w����k����M�ߋ������f����e�0���A�������Y��b��Bq�&Y
��|ڿ+ݒ%g��x��p�@}M��3k�'Z�[��^7��S �1n�m33~�4�ҭ���"{Q6#�&��L��A�j ��z�hP��	E�ǁ�2�z�<�$���@������^ґ|��xp{����<��^��O?�	��\�G�lR�$��Q�,l<�����Ȃ�"df77�'p9��t["@M�H"(�@:3�u�QP�}>%�3G_��k��D|�E�ϫ���dw���9t�H%��_R�����[��/}Ӳ�����/�n���F��8�N ��6Z����.�.U����ȯM/��c�CL�Ӊ �P���U�Bx�JP�7��CF�w�'?�S)-�$'k��/�N�v�Z�J�v9g�����匽[�@�K�ox�t�H�R�c�؆5q<�҆ȳ�jɒ5)��<0[/{�SkB���1�C�ã�n
��{�fⳐ����	�QV|�E����RD*�(��滛��﯏���_z{�),U_Z#��$#"�#^C�!��W�@|����'�S.����~`3��YS�>	�ΘR$~7��q~�����>�(_�������&�a/:�m�;?Q��)��0JPR���$`�y?�W�w=X�8�tz��Zpп�Z��rފ��'�ܧ6���ޭ�q�˧�]�&8	��U��J�\L{`�s�Ue �mO4<�F�����yeo��r︙�������� O+Z7וAHx�Q���d�� �{K����KU{�+�#	"�I~�"B�>�'�'�� ����*P��z=kTw/�m�4Gޞd���,�Zw�G�<��։��8��G"�V7���l�6�̜փ�>�u�]P0�����궠�
*�V�Ftr����BO�h\e��e�zw���r��B�����-g�>Ǖ�e`�<c�	�@���D��)�+9 �EY��/��/��V*#�O�e�#A�4)�1�R����~�8f7a�\�G�g����Y )2��s2��D?Q-�}\���*�QǄ߼�4�7��n��hl�;8�j.ߖA?"����?S��|�r�u�0�0�}���s��L�NR(? h�ߪ���	pOB1a	L	(����]�b*�ĵ��8���y�l��^��B��B�M{��3m��O�rB&_��J;J&��d��Wej���-E�c{���nj��.�n�(>&/f�1;��Mf$�a�c^1�.9o�$#��k�~/1��������<f?k��5'��uD[%�U^��Me�L%��x^�v�ξ�������ѯ��j��"7�7�k�zC\\�&>�&۩'93��bB������=����U�JYu���J@��Z�nEWBވ,�zȥ��4B[�<آ��~��1�t/�K�N�a�I�WS۾&�a�yh�)���G���hYt�����8:/3� #���e/�O&x7�,`;�$הi��,�$�HRa3�rR�2����ᩰ���TJ�����v��#T(=]�x�ȝ(�Ϯ���f����^�pdK?:�	#�i��.7�5m!:II�
�um���7"� ��"�}|�0���gε�q��a	��/��F~��`�i@��*��%�2�v��b�����ݎ$��6���=vW\a���><<�)R���p��Q��43,��A�D�TP�i��(�;�g�	�ȾN��	���=S�E-�M��������	�K'��Re��"Z�<�����(��<�%��z��z�ڸ|A�4�"��ݾw0?~����5٥}�2���d�A�&>ԥ}v��+�����+)�Ǽ�ǚ��i3]�S��Q�i�A2�9י�i�I�2-Ě�b��R�4�a��B�6|���u΍y�Eŗ#��7Ww�L!�ˋ����f��?G�x�ѭu�͠���f�54f0��璨^��1��`U�o}G����}n����d��@u�bix�6���!��e���=�ؗ�uJ�7����)�?��=��*%���l����q~ֿ���n�5�����TXM-�P�m�6?'���佺��ۉ:�B��y�i��T�� k~՚	;�7���b>=�6hZ�yV��o�P��ߘAY�t<q����3�˚�������n�T8�&�GZ���x�d���`���z���"8�\��X2sJo��XR+G�3�I�� 3ؕ��[��V,4����43~�C�j4p�W��u[�@��} j��)�s����e�+*�"��v�Ժ/�
�F�V��D�2������M<��M!��$_!(G!���ݺx%��mM�{��lck� ��m�a>�;�ۛ�4`���=bG�>5Y�=�ʃ��jG���r�o6<�x ���o�s��=�q�ʢC+��Σ{�q�>I�(Sy�H��c�eGM�>�\��g�]��P!(��q-�C�#1�A�%|��A$����AM��7�*��\o�s���0����3��y3�i���7�ww@��47�os;@`2�0�x�k����t+�@%���H��DGI'i�F��|h$�ǝ�j���2D��F>(2{PmqŹ���q]��\:~~�o��ZhF~}�MuF�<����zyP�K6��0�$%����$�^�B�-Jp��eOI�*����%>4cd���#�L��)��-����p�JF�V�Qa�;$�ИW�Zm��d^W��q��)ƭS�0h-�WG��!y����m�	��y��}ܖp5�~�|>�ʿ9N��[U[|��!��XG��,n��O�ˤh/���<�\H����l;Z޻�/�B�#��ˏ$ *7���d/zƝ�Ch�k1��Ӊ�-%��µG�1�p�\�W~ǧ�cpP\ ����䩇/���;���"$T0Y�x��?���
���Ui������� �B�ps��r��ԙ�v��fʂw���? ���g_��[L&	�j���K'��;FbF6Եq9�ތ�h�ĳ ��c�
��#�b&�#t�.�,��C�P�X�U.��5��y�;"0L�<�_��C��tO�So�1^%M&����b��M%��	Ví�G/��W<��yH-�����\�Y��3�=�N��Aw�3��Y��uH?�U��S����ps��Ԓ>�)�����@���F�~����''�@��c�J��$(�k�5���帿'��'Q�%�ǫz�D�U�q��=w��f�v�d��$�Uiiof�»T�$4��loK��]�dX�XN���� BZC�Q&m��=&S�~�#i��(�`@"��*�u����k�;2W>�����qpx�EV��|¾Äua��Eq�V��x)J�p�ߛ|��h"Kh׃�WReS�]��gk��.�ʖ<P��tq�_�d)��`��{Y��|ձO�s5�L��%^!H4��3�x`��*Y��O��x��KT;����%�z���
�t:s�SU)�R.^n�l��@�?���ǧ@	�!���g�|�Z����ԭ��s7�k~�*�q����8��S}�
������R�4»XZς�w�5���A{'f!��YTwK�$%��WTA~�@�m��F%」��ƹ��?�����r#�|�?'DO�y����7�d��ǡp;]%,��C���n��,�LH��܎Y+�$���_����^q���L����\������F<��6��;B���:��5O7��z���x�D�����ìI�t9��A�:@)��,N��O ��UR~$e��r@bz�0�5�d\�mf��H�q�I� ����~�Z�>�.�]t|���F��������p��&�t�#K�Gc��8�P�����9.�D`�<��9�� j�4Q�Y��lw0.F�L�ڗ�ҧ��P���#2[�dX���ه���\q1��7����3�5j�Z�H�!T���O"��f�!%�k����n3ڑ���R���ri1�՚��n��� ���Іra*�v;~���J5�K;�J$,I��VO�b��ݑŀ��P�lA��U:-��H�qh�;M' zw�5M�>���c7�
I�ռ�Z3fmXsir�@��V�]/��ޖ���b`���l��Cڲ�*>Wl�CA�(d����m��W�c̣0<մ�k$א/�!B+���kz5�؂��,9r�eO:0��R]�LqSi�	�o�	|����<��{�Gy�w���7K౑�t2`!�WC��UT֣����P�����,5�+ �:V`57PlE�N`v���ejn"�
�M5��$��Qa�<U�q��0�KV3�S��2]�xi��9��^M���?�Vh�}jV^lZ�(����=��
����a/L���0�Z����e����.���)�yglS����+�~��؍�M��l֧�A�t�Q�/U'H�����s5����V��eՃ�C��ej�a�)��8{�*�o)'ީ��U,]`7t;�qܥ���KtySE�|7���(�%�1[�/~�t���Ż����f�sDHT��-���')���Iu��y��Nh�>���!�y����1$/
'`p��
2�qC��J�&��B�\;�a�*\�~v�	UZ���Ӭ"�N�or�A�pLY�ڠ�`g������Ll��ئ�(�3b�ٳ��9��6w6d�q���9	��E�_�O8#q�2;�Dv��ݜ�9�'��ꨅU�rk.���Bus:�oIs�O��4���	e���>�%�vc������(��x��۵I�8�Ó���n��sI��,#Hf��#E�o���$������&�[��	,�.�Vч:^-T�՛��'���Q|m�o2J�1/���s��F�sh7��Z4;�Vz����11s��oa�:TXs�z{djy�Vk�k	�QD�U�7{������2��v@xC�v��v&��\BQ��|b�+��nr������\�ε�6�Ce#�\�kV��R���k.0�-�M?%�<ӻ��#����
}�MT����:<R(6��6��/Ƭ��c\�k�ɧ%��/�O�� �]�VoZ4_\~�`u�n_L|*�)�U�-4�^\ϻ�#���OT�ҹY4��%!�WF�_>&�zY-Y~�o���1�X���⏜s'`P�<��v�|U!L�C����CF�D��uq�*!)o@4PG�`�]��VmC�n���	U�4K@9t6���*K`?���>3jf�wu��qP$�N���4YHnHG[@�����ۙ�u��a�(�	�R�5�����m̩��1F'���w,�f=v�~o�����v�+g!�o����ON`X�2c�nuȠ���uc&ڰ�C�.�׃�8�7��j���C�r�qb=�������?�S�j�3уɑ�}	���$xrntl鄒�U�	�y�^�<��+,�,(�L_�.+�P��Zm�$]��l��(�3G���`�sC�i�PW���m��S�#<�m�۽B�`(m9q
ûH��k��p��:nr��(�����k]`��SFک�]L��e:��<.�
dis�`���,��7�I
����(%�iS���w��>��[���q�	�^|�1�#��o)��p�E�E�{���i�42��E���)㩱�Ќb�T��ӱ2��Ჿ%���s݄�'�O�KD��q�$�rM�z��22ߜ��&��z诽bPZ�m�R�HdL��Lrc��)������9С�8@j�ֱfW6^+�)�����#�@/�eeT^Γu��h���-1����F�^�M{'�-;<����3�B���� I�y%]%cō�kN�</0�� ����@#�іjԏ�]�@�]j�}�$����|T-�.}(`��Tx�k�{·�ѱF�V�b�Y� ���"���,)���}�HI���)�q�z�����ٖ.�/���������[���w��I4�����d�,ZG7�X��5�n��-�q��I�	hH�s���P�f�h[@�G�G-|��kU4%E�~{����G7|�)ű���ݥ)�If�YBH��Usz�S�u�/a�Ջ��Q�����Ȟ=2��i�5���?�a}O���R�s�)��m��v�S�&��L4���[���ItY2	��g�	�k�b�ut3��+�T}�M&g�π�C��
����֥��s���0�y�3��J�����ڕ�#t1D���_���M�h�>�X�f�3������e� �R^�n�����g��ۍ�{�����k�>��Woc����F�U��X�
z[�ntnKN�J�1H�Ř�� {�g��B[)p�
�&~k�ldd?(���6*?��k��}�a1��^�DN4������*�2m%5g2m��2�\(A������8��aB��|Ĥp�Y���q��+�֫���m���I��v���h&б��x�3�N:7^�@�/��@��-�pYa?�^�����2TC�;��V9�RI�7s�ˍƖ�B���5h��n����:sq*�O�{�P���J����!�)D٘r%q�0�MG\%8�}�c5u��~�0������|"��.�+� �^'���ɑ�z�Ȥ؄�t����OT�	��弡_'�ѣ�[CF��3���8���-��Kl���VV�ٌAE���T08
�Fi�4Op��@��pf��{�<��p��37}j�@.��:�W�7���qBr���h�֯:dM(�AP�Ut�T}��Jyl�V:�����D2�䵥��Yx���A�KfZ���� /Q����׫ו� s�x�\����3���>��[MPL��B*����,"��g<��'\P���[���x�w�2�5M�2e4���I����|F�|]賷D+ذ���0.2y �gU:& ���������JH��*�J\1}n����� �qɔ�R�Y
�=�$yd
(�z�`g�('����3"����L�7
B�M�%A{4�`H�;��Yf��=��rP-��G����v�CRM`��5�B�[���urZQ�%�]��� �)/~��~k{��Ez̐�e��o�!(^����6���C�dY�H�o;��\U��P�w�s[�zt��X�F�2b,�x.s�S2-�-P�_M"��25����dD�Q�zT�=~9[���2��W0:�ϐ-)V�	~T+��U&�1�=�ѐ�㈿C�؅t9���QPOR@}�m�ܿ�c!aC�>�B7LϦ